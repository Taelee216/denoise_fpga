

module gru2( noise_gru_state, noise_input, clk );

	parameter 			float = 32;

	reg		[          float : 0]	noise_gru_bias_array[143:0];
	wire	[(  144*float)-1 : 0]	noise_gru_bias;

	reg		[          float : 0]	noise_gru_input_weights_array[12959:0];
	wire	[(12960*float)-1 : 0]	noise_gru_input_weights;

	reg		[          float : 0]	noise_gru_recurrent_weights_array[6911:0];
	wire	[( 6912*float)-1 : 0]	noise_gru_recurrent_weights;


	output 	[(   48*float)-1 : 0]	noise_gru_state;
	input 	[(   90*float)-1 : 0]	noise_input;
	input 				clk;

	
	reg 	[(   90*float)-1 : 0]	z ,tmpz, r, tmpr, h, tmph, tmptmp;

	reg		[        float-1 : 0]	weights_scale;
	reg		[(   48*float)-1 : 0]	sum, tmpsum1, tmpsum2;

	integer	index1		= 0;
	integer	index2		= 0;
	integer	index3		= 0;
	integer	M		= 90;
	integer	N		= 48;
	integer	stride		= 144;
	integer	one		= 1;

/////////////////////////////////////////////////////////////////////////////////////////////////////
{
	assign	noise_gru_bias_array[    0] = 32'b01000010010011000000000000000000;
	assign	noise_gru_bias_array[    1] = 32'b01000010000000000000000000000000;
	assign	noise_gru_bias_array[    2] = 32'b01000010101100000000000000000000;
	assign	noise_gru_bias_array[    3] = 32'b01000010011100000000000000000000;
	assign	noise_gru_bias_array[    4] = 32'b11000010100000000000000000000000;
	assign	noise_gru_bias_array[    5] = 32'b01000010101110000000000000000000;
	assign	noise_gru_bias_array[    6] = 32'b01000000101000000000000000000000;
	assign	noise_gru_bias_array[    7] = 32'b11000010000100000000000000000000;
	assign	noise_gru_bias_array[    8] = 32'b11000010010001000000000000000000;
	assign	noise_gru_bias_array[    9] = 32'b01000010101111100000000000000000;
	assign	noise_gru_bias_array[   10] = 32'b01000010110011000000000000000000;
	assign	noise_gru_bias_array[   11] = 32'b11000001101000000000000000000000;
	assign	noise_gru_bias_array[   12] = 32'b10111111100000000000000000000000;
	assign	noise_gru_bias_array[   13] = 32'b01000001011000000000000000000000;
	assign	noise_gru_bias_array[   14] = 32'b01000001000000000000000000000000;
	assign	noise_gru_bias_array[   15] = 32'b01000001101010000000000000000000;
	assign	noise_gru_bias_array[   16] = 32'b11000010000100000000000000000000;
	assign	noise_gru_bias_array[   17] = 32'b11000010100010000000000000000000;
	assign	noise_gru_bias_array[   18] = 32'b01000010011110000000000000000000;
	assign	noise_gru_bias_array[   19] = 32'b01000010001110000000000000000000;
	assign	noise_gru_bias_array[   20] = 32'b01000001001000000000000000000000;
	assign	noise_gru_bias_array[   21] = 32'b11000010011100000000000000000000;
	assign	noise_gru_bias_array[   22] = 32'b11000010110011100000000000000000;
	assign	noise_gru_bias_array[   23] = 32'b11000001100000000000000000000000;
	assign	noise_gru_bias_array[   24] = 32'b11000001111100000000000000000000;
	assign	noise_gru_bias_array[   25] = 32'b11000010001010000000000000000000;
	assign	noise_gru_bias_array[   26] = 32'b11000010001011000000000000000000;
	assign	noise_gru_bias_array[   27] = 32'b01000010000011000000000000000000;
	assign	noise_gru_bias_array[   28] = 32'b11000000100000000000000000000000;
	assign	noise_gru_bias_array[   29] = 32'b01000001101110000000000000000000;
	assign	noise_gru_bias_array[   30] = 32'b01000010110000100000000000000000;
	assign	noise_gru_bias_array[   31] = 32'b01000010001110000000000000000000;
	assign	noise_gru_bias_array[   32] = 32'b11000001111010000000000000000000;
	assign	noise_gru_bias_array[   33] = 32'b11000001100000000000000000000000;
	assign	noise_gru_bias_array[   34] = 32'b01000010100011100000000000000000;
	assign	noise_gru_bias_array[   35] = 32'b01000010010100000000000000000000;
	assign	noise_gru_bias_array[   36] = 32'b11000001101000000000000000000000;
	assign	noise_gru_bias_array[   37] = 32'b11000001101110000000000000000000;
	assign	noise_gru_bias_array[   38] = 32'b01000010101101100000000000000000;
	assign	noise_gru_bias_array[   39] = 32'b01000001100000000000000000000000;
	assign	noise_gru_bias_array[   40] = 32'b01000010100010100000000000000000;
	assign	noise_gru_bias_array[   41] = 32'b11000001010100000000000000000000;
	assign	noise_gru_bias_array[   42] = 32'b11000001101110000000000000000000;
	assign	noise_gru_bias_array[   43] = 32'b01000010100100100000000000000000;
	assign	noise_gru_bias_array[   44] = 32'b11000001100010000000000000000000;
	assign	noise_gru_bias_array[   45] = 32'b01000001010100000000000000000000;
	assign	noise_gru_bias_array[   46] = 32'b01000001111100000000000000000000;
	assign	noise_gru_bias_array[   47] = 32'b01000001101110000000000000000000;
	assign	noise_gru_bias_array[   48] = 32'b00111111100000000000000000000000;
	assign	noise_gru_bias_array[   49] = 32'b11000001110110000000000000000000;
	assign	noise_gru_bias_array[   50] = 32'b01000010010101000000000000000000;
	assign	noise_gru_bias_array[   51] = 32'b11000001110000000000000000000000;
	assign	noise_gru_bias_array[   52] = 32'b11000010100011100000000000000000;
	assign	noise_gru_bias_array[   53] = 32'b01000010001101000000000000000000;
	assign	noise_gru_bias_array[   54] = 32'b01000010001010000000000000000000;
	assign	noise_gru_bias_array[   55] = 32'b11000010010001000000000000000000;
	assign	noise_gru_bias_array[   56] = 32'b01000001111000000000000000000000;
	assign	noise_gru_bias_array[   57] = 32'b11000001100000000000000000000000;
	assign	noise_gru_bias_array[   58] = 32'b11000001101000000000000000000000;
	assign	noise_gru_bias_array[   59] = 32'b01000010011101000000000000000000;
	assign	noise_gru_bias_array[   60] = 32'b01000010001000000000000000000000;
	assign	noise_gru_bias_array[   61] = 32'b11000010110100000000000000000000;
	assign	noise_gru_bias_array[   62] = 32'b01000010010110000000000000000000;
	assign	noise_gru_bias_array[   63] = 32'b11000000101000000000000000000000;
	assign	noise_gru_bias_array[   64] = 32'b01000001111110000000000000000000;
	assign	noise_gru_bias_array[   65] = 32'b01000001001000000000000000000000;
	assign	noise_gru_bias_array[   66] = 32'b11000010010011000000000000000000;
	assign	noise_gru_bias_array[   67] = 32'b11000010000101000000000000000000;
	assign	noise_gru_bias_array[   68] = 32'b11000000110000000000000000000000;
	assign	noise_gru_bias_array[   69] = 32'b11000010101010100000000000000000;
	assign	noise_gru_bias_array[   70] = 32'b01000001000100000000000000000000;
	assign	noise_gru_bias_array[   71] = 32'b01000010010011000000000000000000;
	assign	noise_gru_bias_array[   72] = 32'b01000001100000000000000000000000;
	assign	noise_gru_bias_array[   73] = 32'b01000000000000000000000000000000;
	assign	noise_gru_bias_array[   74] = 32'b11000001110100000000000000000000;
	assign	noise_gru_bias_array[   75] = 32'b01000010011000000000000000000000;
	assign	noise_gru_bias_array[   76] = 32'b11000010000111000000000000000000;
	assign	noise_gru_bias_array[   77] = 32'b11000000101000000000000000000000;
	assign	noise_gru_bias_array[   78] = 32'b11000001110110000000000000000000;
	assign	noise_gru_bias_array[   79] = 32'b11000001010100000000000000000000;
	assign	noise_gru_bias_array[   80] = 32'b11000010010001000000000000000000;
	assign	noise_gru_bias_array[   81] = 32'b01000001111100000000000000000000;
	assign	noise_gru_bias_array[   82] = 32'b01000000100000000000000000000000;
	assign	noise_gru_bias_array[   83] = 32'b11000010100000000000000000000000;
	assign	noise_gru_bias_array[   84] = 32'b11000010001001000000000000000000;
	assign	noise_gru_bias_array[   85] = 32'b01000010001101000000000000000000;
	assign	noise_gru_bias_array[   86] = 32'b11000001101110000000000000000000;
	assign	noise_gru_bias_array[   87] = 32'b01000001011000000000000000000000;
	assign	noise_gru_bias_array[   88] = 32'b11000001100110000000000000000000;
	assign	noise_gru_bias_array[   89] = 32'b11000001001000000000000000000000;
	assign	noise_gru_bias_array[   90] = 32'b11000010010111000000000000000000;
	assign	noise_gru_bias_array[   91] = 32'b11000010011101000000000000000000;
	assign	noise_gru_bias_array[   92] = 32'b11000010000011000000000000000000;
	assign	noise_gru_bias_array[   93] = 32'b01000010001110000000000000000000;
	assign	noise_gru_bias_array[   94] = 32'b11000001111110000000000000000000;
	assign	noise_gru_bias_array[   95] = 32'b11000001010000000000000000000000;
	assign	noise_gru_bias_array[   96] = 32'b11000010101110100000000000000000;
	assign	noise_gru_bias_array[   97] = 32'b11000001111000000000000000000000;
	assign	noise_gru_bias_array[   98] = 32'b01000001001100000000000000000000;
	assign	noise_gru_bias_array[   99] = 32'b11000000110000000000000000000000;
	assign	noise_gru_bias_array[  100] = 32'b11000010001110000000000000000000;
	assign	noise_gru_bias_array[  101] = 32'b11000001010000000000000000000000;
	assign	noise_gru_bias_array[  102] = 32'b00111111100000000000000000000000;
	assign	noise_gru_bias_array[  103] = 32'b01000001011100000000000000000000;
	assign	noise_gru_bias_array[  104] = 32'b11000010000101000000000000000000;
	assign	noise_gru_bias_array[  105] = 32'b11000010110101100000000000000000;
	assign	noise_gru_bias_array[  106] = 32'b11000010010010000000000000000000;
	assign	noise_gru_bias_array[  107] = 32'b01000000010000000000000000000000;
	assign	noise_gru_bias_array[  108] = 32'b01000010010110000000000000000000;
	assign	noise_gru_bias_array[  109] = 32'b11000001110100000000000000000000;
	assign	noise_gru_bias_array[  110] = 32'b11000010101011000000000000000000;
	assign	noise_gru_bias_array[  111] = 32'b01000001011000000000000000000000;
	assign	noise_gru_bias_array[  112] = 32'b01000010100001000000000000000000;
	assign	noise_gru_bias_array[  113] = 32'b11000010010110000000000000000000;
	assign	noise_gru_bias_array[  114] = 32'b11000010000110000000000000000000;
	assign	noise_gru_bias_array[  115] = 32'b11000010100011000000000000000000;
	assign	noise_gru_bias_array[  116] = 32'b10111111100000000000000000000000;
	assign	noise_gru_bias_array[  117] = 32'b01000010100010100000000000000000;
	assign	noise_gru_bias_array[  118] = 32'b01000010001110000000000000000000;
	assign	noise_gru_bias_array[  119] = 32'b11000001010000000000000000000000;
	assign	noise_gru_bias_array[  120] = 32'b11000011000000000000000000000000;
	assign	noise_gru_bias_array[  121] = 32'b11000010010111000000000000000000;
	assign	noise_gru_bias_array[  122] = 32'b00000000000000000000000000000000;
	assign	noise_gru_bias_array[  123] = 32'b01000001100010000000000000000000;
	assign	noise_gru_bias_array[  124] = 32'b01000010010000000000000000000000;
	assign	noise_gru_bias_array[  125] = 32'b11000010100000000000000000000000;
	assign	noise_gru_bias_array[  126] = 32'b11000001110000000000000000000000;
	assign	noise_gru_bias_array[  127] = 32'b01000001000100000000000000000000;
	assign	noise_gru_bias_array[  128] = 32'b11000010100001100000000000000000;
	assign	noise_gru_bias_array[  129] = 32'b11000010110101100000000000000000;
	assign	noise_gru_bias_array[  130] = 32'b11000010110010100000000000000000;
	assign	noise_gru_bias_array[  131] = 32'b11000010001011000000000000000000;
	assign	noise_gru_bias_array[  132] = 32'b11000000100000000000000000000000;
	assign	noise_gru_bias_array[  133] = 32'b01000010101000000000000000000000;
	assign	noise_gru_bias_array[  134] = 32'b11000010010100000000000000000000;
	assign	noise_gru_bias_array[  135] = 32'b11000010101101000000000000000000;
	assign	noise_gru_bias_array[  136] = 32'b11000001101110000000000000000000;
	assign	noise_gru_bias_array[  137] = 32'b11000010100000000000000000000000;
	assign	noise_gru_bias_array[  138] = 32'b01000001111110000000000000000000;
	assign	noise_gru_bias_array[  139] = 32'b01000010101011000000000000000000;
	assign	noise_gru_bias_array[  140] = 32'b11000010010010000000000000000000;
	assign	noise_gru_bias_array[  141] = 32'b01000000000000000000000000000000;
	assign	noise_gru_bias_array[  142] = 32'b11000010000110000000000000000000;
	assign	noise_gru_bias_array[  143] = 32'b01000000111000000000000000000000;

	assign	noise_gru_input_weights_array[    0] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[    1] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[    2] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[    3] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[    4] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[    5] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[    6] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[    7] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[    8] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[    9] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[   10] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[   11] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[   12] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[   13] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[   14] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[   15] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[   16] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[   17] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[   18] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[   19] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[   20] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[   21] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[   22] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[   23] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[   24] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[   25] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[   26] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[   27] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[   28] = 32'b01000010111000000000000000000000;
	assign	noise_gru_input_weights_array[   29] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[   30] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[   31] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[   32] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[   33] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[   34] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[   35] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[   36] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[   37] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[   38] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[   39] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[   40] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[   41] = 32'b11000010110001100000000000000000;
	assign	noise_gru_input_weights_array[   42] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[   43] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[   44] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[   45] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[   46] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[   47] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[   48] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[   49] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[   50] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[   51] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[   52] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[   53] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[   54] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[   55] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[   56] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[   57] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[   58] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[   59] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[   60] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[   61] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[   62] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[   63] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[   64] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[   65] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[   66] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[   67] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[   68] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[   69] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[   70] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[   71] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[   72] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[   73] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[   74] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[   75] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[   76] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[   77] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[   78] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[   79] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[   80] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[   81] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[   82] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[   83] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[   84] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[   85] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[   86] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[   87] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[   88] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[   89] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[   90] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[   91] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[   92] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[   93] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[   94] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[   95] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[   96] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[   97] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[   98] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[   99] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[  100] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[  101] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[  102] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[  103] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[  104] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[  105] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[  106] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[  107] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[  108] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[  109] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[  110] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[  111] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[  112] = 32'b01000010110100000000000000000000;
	assign	noise_gru_input_weights_array[  113] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[  114] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[  115] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[  116] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[  117] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[  118] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[  119] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[  120] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[  121] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[  122] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[  123] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[  124] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[  125] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[  126] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[  127] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[  128] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[  129] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[  130] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[  131] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[  132] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[  133] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[  134] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[  135] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[  136] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[  137] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[  138] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[  139] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[  140] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[  141] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[  142] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[  143] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[  144] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[  145] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[  146] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[  147] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[  148] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[  149] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[  150] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[  151] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[  152] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[  153] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[  154] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[  155] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[  156] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[  157] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[  158] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[  159] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[  160] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[  161] = 32'b11000010110111000000000000000000;
	assign	noise_gru_input_weights_array[  162] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[  163] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[  164] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[  165] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[  166] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[  167] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[  168] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[  169] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[  170] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[  171] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[  172] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[  173] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[  174] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[  175] = 32'b11000010111001000000000000000000;
	assign	noise_gru_input_weights_array[  176] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[  177] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[  178] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[  179] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[  180] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[  181] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[  182] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[  183] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[  184] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[  185] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[  186] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[  187] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[  188] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[  189] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[  190] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[  191] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[  192] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[  193] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[  194] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[  195] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[  196] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[  197] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[  198] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[  199] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[  200] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[  201] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[  202] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[  203] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[  204] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[  205] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[  206] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[  207] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[  208] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[  209] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[  210] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[  211] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[  212] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[  213] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[  214] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[  215] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[  216] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[  217] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[  218] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[  219] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[  220] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[  221] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[  222] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[  223] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[  224] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[  225] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[  226] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[  227] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[  228] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[  229] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[  230] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[  231] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[  232] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[  233] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[  234] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[  235] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[  236] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[  237] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[  238] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[  239] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[  240] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[  241] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[  242] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[  243] = 32'b11000010110101000000000000000000;
	assign	noise_gru_input_weights_array[  244] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[  245] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[  246] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[  247] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[  248] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[  249] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[  250] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[  251] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[  252] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[  253] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[  254] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[  255] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[  256] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[  257] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[  258] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[  259] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[  260] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[  261] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[  262] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[  263] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[  264] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[  265] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[  266] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[  267] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[  268] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[  269] = 32'b11000010110110000000000000000000;
	assign	noise_gru_input_weights_array[  270] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[  271] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[  272] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[  273] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[  274] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[  275] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[  276] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[  277] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[  278] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[  279] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[  280] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[  281] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[  282] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[  283] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[  284] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[  285] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[  286] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[  287] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[  288] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[  289] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[  290] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[  291] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[  292] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[  293] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[  294] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[  295] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[  296] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[  297] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[  298] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[  299] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[  300] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[  301] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[  302] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[  303] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[  304] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[  305] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[  306] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[  307] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[  308] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[  309] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[  310] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[  311] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[  312] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[  313] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[  314] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[  315] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[  316] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[  317] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[  318] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[  319] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[  320] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[  321] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[  322] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[  323] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[  324] = 32'b01000010110100100000000000000000;
	assign	noise_gru_input_weights_array[  325] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[  326] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[  327] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[  328] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[  329] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[  330] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[  331] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[  332] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[  333] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[  334] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[  335] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[  336] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[  337] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[  338] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[  339] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[  340] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[  341] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[  342] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[  343] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[  344] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[  345] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[  346] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[  347] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[  348] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[  349] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[  350] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[  351] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[  352] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[  353] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[  354] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[  355] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[  356] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[  357] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[  358] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[  359] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[  360] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[  361] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[  362] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[  363] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[  364] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[  365] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[  366] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[  367] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[  368] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[  369] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[  370] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[  371] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[  372] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[  373] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[  374] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[  375] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[  376] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[  377] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[  378] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[  379] = 32'b11000010101110000000000000000000;
	assign	noise_gru_input_weights_array[  380] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[  381] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[  382] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[  383] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[  384] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[  385] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[  386] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[  387] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[  388] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[  389] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[  390] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[  391] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[  392] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[  393] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[  394] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[  395] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[  396] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[  397] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[  398] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[  399] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[  400] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[  401] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[  402] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[  403] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[  404] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[  405] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[  406] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[  407] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[  408] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[  409] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[  410] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[  411] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[  412] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[  413] = 32'b11000010110010100000000000000000;
	assign	noise_gru_input_weights_array[  414] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[  415] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[  416] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[  417] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[  418] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[  419] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[  420] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[  421] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[  422] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[  423] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[  424] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[  425] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[  426] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[  427] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[  428] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[  429] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[  430] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[  431] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[  432] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[  433] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[  434] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[  435] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[  436] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[  437] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[  438] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[  439] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[  440] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[  441] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[  442] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[  443] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[  444] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[  445] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[  446] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[  447] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[  448] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[  449] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[  450] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[  451] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[  452] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[  453] = 32'b11000010110111100000000000000000;
	assign	noise_gru_input_weights_array[  454] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[  455] = 32'b11000010101110000000000000000000;
	assign	noise_gru_input_weights_array[  456] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[  457] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[  458] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[  459] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[  460] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[  461] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[  462] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[  463] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[  464] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[  465] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[  466] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[  467] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[  468] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[  469] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[  470] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[  471] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[  472] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[  473] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[  474] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[  475] = 32'b11000010110110100000000000000000;
	assign	noise_gru_input_weights_array[  476] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[  477] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[  478] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[  479] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[  480] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[  481] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[  482] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[  483] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[  484] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[  485] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[  486] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[  487] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[  488] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[  489] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[  490] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[  491] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[  492] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[  493] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[  494] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[  495] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[  496] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[  497] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[  498] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[  499] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[  500] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[  501] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[  502] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[  503] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[  504] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[  505] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[  506] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[  507] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[  508] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[  509] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[  510] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[  511] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[  512] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[  513] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[  514] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[  515] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[  516] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[  517] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[  518] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[  519] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[  520] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[  521] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[  522] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[  523] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[  524] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[  525] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[  526] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[  527] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[  528] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[  529] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[  530] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[  531] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[  532] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[  533] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[  534] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[  535] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[  536] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[  537] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[  538] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[  539] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[  540] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[  541] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[  542] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[  543] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[  544] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[  545] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[  546] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[  547] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[  548] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[  549] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[  550] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[  551] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[  552] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[  553] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[  554] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[  555] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[  556] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[  557] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[  558] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[  559] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[  560] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[  561] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[  562] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[  563] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[  564] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[  565] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[  566] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[  567] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[  568] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[  569] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[  570] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[  571] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[  572] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[  573] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[  574] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[  575] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[  576] = 32'b01000010101111000000000000000000;
	assign	noise_gru_input_weights_array[  577] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[  578] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[  579] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[  580] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[  581] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[  582] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[  583] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[  584] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[  585] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[  586] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[  587] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[  588] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[  589] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[  590] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[  591] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[  592] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[  593] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[  594] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[  595] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[  596] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[  597] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[  598] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[  599] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[  600] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[  601] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[  602] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[  603] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[  604] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[  605] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[  606] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[  607] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[  608] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[  609] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[  610] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[  611] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[  612] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[  613] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[  614] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[  615] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[  616] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[  617] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[  618] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[  619] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[  620] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[  621] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[  622] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[  623] = 32'b01000010110000000000000000000000;
	assign	noise_gru_input_weights_array[  624] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[  625] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[  626] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[  627] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[  628] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[  629] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[  630] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[  631] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[  632] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[  633] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[  634] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[  635] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[  636] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[  637] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[  638] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[  639] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[  640] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[  641] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[  642] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[  643] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[  644] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[  645] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[  646] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[  647] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[  648] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[  649] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[  650] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[  651] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[  652] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[  653] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[  654] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[  655] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[  656] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[  657] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[  658] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[  659] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[  660] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[  661] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[  662] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[  663] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[  664] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[  665] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[  666] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[  667] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[  668] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[  669] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[  670] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[  671] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[  672] = 32'b11000010110011000000000000000000;
	assign	noise_gru_input_weights_array[  673] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[  674] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[  675] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[  676] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[  677] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[  678] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[  679] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[  680] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[  681] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[  682] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[  683] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[  684] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[  685] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[  686] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[  687] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[  688] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[  689] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[  690] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[  691] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[  692] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[  693] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[  694] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[  695] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[  696] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[  697] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[  698] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[  699] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[  700] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[  701] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[  702] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[  703] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[  704] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[  705] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[  706] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[  707] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[  708] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[  709] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[  710] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[  711] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[  712] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[  713] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[  714] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[  715] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[  716] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[  717] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[  718] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[  719] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[  720] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[  721] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[  722] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[  723] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[  724] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[  725] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[  726] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[  727] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[  728] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[  729] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[  730] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[  731] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[  732] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[  733] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[  734] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[  735] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[  736] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[  737] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[  738] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[  739] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[  740] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[  741] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[  742] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[  743] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[  744] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[  745] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[  746] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[  747] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[  748] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[  749] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[  750] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[  751] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[  752] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[  753] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[  754] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[  755] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[  756] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[  757] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[  758] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[  759] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[  760] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[  761] = 32'b01000010110010000000000000000000;
	assign	noise_gru_input_weights_array[  762] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[  763] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[  764] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[  765] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[  766] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[  767] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[  768] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[  769] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[  770] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[  771] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[  772] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[  773] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[  774] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[  775] = 32'b01000010101111000000000000000000;
	assign	noise_gru_input_weights_array[  776] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[  777] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[  778] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[  779] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[  780] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[  781] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[  782] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[  783] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[  784] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[  785] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[  786] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[  787] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[  788] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[  789] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[  790] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[  791] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[  792] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[  793] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[  794] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[  795] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[  796] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[  797] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[  798] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[  799] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[  800] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[  801] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[  802] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[  803] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[  804] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[  805] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[  806] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[  807] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[  808] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[  809] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[  810] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[  811] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[  812] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[  813] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[  814] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[  815] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[  816] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[  817] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[  818] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[  819] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[  820] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[  821] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[  822] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[  823] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[  824] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[  825] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[  826] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[  827] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[  828] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[  829] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[  830] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[  831] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[  832] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[  833] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[  834] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[  835] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[  836] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[  837] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[  838] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[  839] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[  840] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[  841] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[  842] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[  843] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[  844] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[  845] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[  846] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[  847] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[  848] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[  849] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[  850] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[  851] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[  852] = 32'b11000010110010100000000000000000;
	assign	noise_gru_input_weights_array[  853] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[  854] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[  855] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[  856] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[  857] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[  858] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[  859] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[  860] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[  861] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[  862] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[  863] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[  864] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[  865] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[  866] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[  867] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[  868] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[  869] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[  870] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[  871] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[  872] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[  873] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[  874] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[  875] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[  876] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[  877] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[  878] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[  879] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[  880] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[  881] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[  882] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[  883] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[  884] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[  885] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[  886] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[  887] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[  888] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[  889] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[  890] = 32'b01000010110100100000000000000000;
	assign	noise_gru_input_weights_array[  891] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[  892] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[  893] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[  894] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[  895] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[  896] = 32'b11000010110001100000000000000000;
	assign	noise_gru_input_weights_array[  897] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[  898] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[  899] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[  900] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[  901] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[  902] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[  903] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[  904] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[  905] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[  906] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[  907] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[  908] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[  909] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[  910] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[  911] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[  912] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[  913] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[  914] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[  915] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[  916] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[  917] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[  918] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[  919] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[  920] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[  921] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[  922] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[  923] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[  924] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[  925] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[  926] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[  927] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[  928] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[  929] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[  930] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[  931] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[  932] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[  933] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[  934] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[  935] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[  936] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[  937] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[  938] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[  939] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[  940] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[  941] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[  942] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[  943] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[  944] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[  945] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[  946] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[  947] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[  948] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[  949] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[  950] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[  951] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[  952] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[  953] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[  954] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[  955] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[  956] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[  957] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[  958] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[  959] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[  960] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[  961] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[  962] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[  963] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[  964] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[  965] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[  966] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[  967] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[  968] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[  969] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[  970] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[  971] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[  972] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[  973] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[  974] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[  975] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[  976] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[  977] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[  978] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[  979] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[  980] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[  981] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[  982] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[  983] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[  984] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[  985] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[  986] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[  987] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[  988] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[  989] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[  990] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[  991] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[  992] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[  993] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[  994] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[  995] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[  996] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[  997] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[  998] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[  999] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 1000] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1001] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1002] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 1003] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 1004] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1005] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1006] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1007] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1008] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 1009] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1010] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 1011] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1012] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1013] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 1014] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1015] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1016] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 1017] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1018] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1019] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1020] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1021] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 1022] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 1023] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 1024] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 1025] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 1026] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 1027] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 1028] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1029] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 1030] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1031] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1032] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1033] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1034] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 1035] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 1036] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 1037] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1038] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1039] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 1040] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 1041] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1042] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 1043] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 1044] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1045] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 1046] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1047] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 1048] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1049] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1050] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 1051] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 1052] = 32'b01000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 1053] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 1054] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 1055] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 1056] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1057] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 1058] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1059] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1060] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 1061] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1062] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1063] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 1064] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 1065] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1066] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1067] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1068] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 1069] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 1070] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1071] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1072] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 1073] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1074] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1075] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 1076] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1077] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 1078] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1079] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 1080] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 1081] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1082] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 1083] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 1084] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 1085] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1086] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1087] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 1088] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 1089] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1090] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 1091] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 1092] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1093] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1094] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1095] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1096] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1097] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 1098] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 1099] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 1100] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 1101] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[ 1102] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 1103] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 1104] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 1105] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1106] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 1107] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 1108] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1109] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 1110] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 1111] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1112] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 1113] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1114] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 1115] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1116] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1117] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1118] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 1119] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 1120] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1121] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 1122] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1123] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1124] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1125] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 1126] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 1127] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1128] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[ 1129] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1130] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1131] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1132] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1133] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1134] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 1135] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1136] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1137] = 32'b01000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1138] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1139] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1140] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 1141] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1142] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1143] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 1144] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1145] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1146] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 1147] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 1148] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 1149] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 1150] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 1151] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 1152] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 1153] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 1154] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 1155] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 1156] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 1157] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 1158] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1159] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 1160] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1161] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 1162] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 1163] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1164] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 1165] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 1166] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1167] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1168] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 1169] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 1170] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 1171] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 1172] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 1173] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1174] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1175] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 1176] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1177] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 1178] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 1179] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1180] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 1181] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1182] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 1183] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1184] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1185] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 1186] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 1187] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1188] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 1189] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 1190] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 1191] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1192] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 1193] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 1194] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1195] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 1196] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 1197] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 1198] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 1199] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1200] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1201] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 1202] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1203] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1204] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 1205] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1206] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1207] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1208] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 1209] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 1210] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 1211] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1212] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 1213] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1214] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 1215] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1216] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 1217] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 1218] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1219] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1220] = 32'b11000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 1221] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 1222] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 1223] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 1224] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1225] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1226] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 1227] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 1228] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 1229] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1230] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1231] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 1232] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 1233] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1234] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 1235] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1236] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 1237] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 1238] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 1239] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 1240] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 1241] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1242] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1243] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 1244] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 1245] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 1246] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1247] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 1248] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1249] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 1250] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1251] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1252] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 1253] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 1254] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1255] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 1256] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1257] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1258] = 32'b11000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 1259] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 1260] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1261] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 1262] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1263] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 1264] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 1265] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 1266] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 1267] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 1268] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1269] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1270] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1271] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1272] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1273] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 1274] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 1275] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 1276] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1277] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 1278] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1279] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1280] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1281] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1282] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 1283] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 1284] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 1285] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 1286] = 32'b11000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 1287] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1288] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1289] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 1290] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1291] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 1292] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 1293] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1294] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 1295] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 1296] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1297] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 1298] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1299] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 1300] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 1301] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1302] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 1303] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 1304] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 1305] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 1306] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 1307] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 1308] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 1309] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 1310] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 1311] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1312] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 1313] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1314] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1315] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1316] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 1317] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 1318] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1319] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1320] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 1321] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 1322] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 1323] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 1324] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1325] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 1326] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1327] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 1328] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 1329] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1330] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 1331] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1332] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1333] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1334] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 1335] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1336] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 1337] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 1338] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 1339] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 1340] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 1341] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 1342] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 1343] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1344] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1345] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 1346] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 1347] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 1348] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 1349] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 1350] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1351] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 1352] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 1353] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 1354] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 1355] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1356] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1357] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 1358] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 1359] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 1360] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 1361] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1362] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1363] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 1364] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 1365] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1366] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1367] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1368] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1369] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 1370] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1371] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1372] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1373] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1374] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 1375] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 1376] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1377] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1378] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 1379] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 1380] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 1381] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1382] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1383] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1384] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 1385] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1386] = 32'b01000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 1387] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 1388] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1389] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 1390] = 32'b01000010110111000000000000000000;
	assign	noise_gru_input_weights_array[ 1391] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 1392] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 1393] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1394] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 1395] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1396] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 1397] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 1398] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 1399] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 1400] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 1401] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1402] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1403] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 1404] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 1405] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 1406] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1407] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1408] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 1409] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1410] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1411] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1412] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 1413] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1414] = 32'b11000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 1415] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 1416] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 1417] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 1418] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1419] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 1420] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 1421] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1422] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1423] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 1424] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1425] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1426] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 1427] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1428] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1429] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 1430] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 1431] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 1432] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1433] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 1434] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 1435] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 1436] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 1437] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1438] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 1439] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 1440] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 1441] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 1442] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1443] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 1444] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1445] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 1446] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 1447] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1448] = 32'b11000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 1449] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 1450] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 1451] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1452] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 1453] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1454] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 1455] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 1456] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 1457] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 1458] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 1459] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 1460] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 1461] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1462] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 1463] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1464] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1465] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1466] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1467] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 1468] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 1469] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1470] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 1471] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 1472] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 1473] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 1474] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1475] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 1476] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1477] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1478] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 1479] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1480] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1481] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 1482] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 1483] = 32'b11000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 1484] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 1485] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 1486] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1487] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 1488] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 1489] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 1490] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 1491] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1492] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 1493] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1494] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 1495] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 1496] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1497] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1498] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 1499] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1500] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 1501] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 1502] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 1503] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1504] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 1505] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1506] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 1507] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1508] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 1509] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 1510] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 1511] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1512] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1513] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 1514] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1515] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 1516] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 1517] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 1518] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1519] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 1520] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1521] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1522] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 1523] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 1524] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 1525] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 1526] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 1527] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 1528] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1529] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1530] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1531] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 1532] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1533] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1534] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 1535] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1536] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 1537] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 1538] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 1539] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1540] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 1541] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 1542] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 1543] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 1544] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 1545] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 1546] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1547] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 1548] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1549] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 1550] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1551] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1552] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1553] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 1554] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1555] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1556] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 1557] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1558] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1559] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1560] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 1561] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 1562] = 32'b01000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 1563] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 1564] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 1565] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1566] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1567] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 1568] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 1569] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 1570] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1571] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 1572] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 1573] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 1574] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 1575] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 1576] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1577] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 1578] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1579] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1580] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1581] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1582] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 1583] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 1584] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1585] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 1586] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1587] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 1588] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 1589] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 1590] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1591] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 1592] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 1593] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 1594] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 1595] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 1596] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1597] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 1598] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 1599] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1600] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1601] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 1602] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 1603] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 1604] = 32'b11000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 1605] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 1606] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 1607] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 1608] = 32'b01000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 1609] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 1610] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 1611] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 1612] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1613] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1614] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 1615] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1616] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 1617] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 1618] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 1619] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 1620] = 32'b01000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 1621] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1622] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1623] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 1624] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1625] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1626] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 1627] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 1628] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1629] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1630] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 1631] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1632] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 1633] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 1634] = 32'b11000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 1635] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1636] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 1637] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1638] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 1639] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 1640] = 32'b01000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 1641] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1642] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 1643] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 1644] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 1645] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1646] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 1647] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1648] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 1649] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 1650] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 1651] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 1652] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1653] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 1654] = 32'b11000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 1655] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 1656] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 1657] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 1658] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 1659] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1660] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 1661] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 1662] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 1663] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1664] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 1665] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 1666] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1667] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1668] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1669] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1670] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1671] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 1672] = 32'b11000010110010100000000000000000;
	assign	noise_gru_input_weights_array[ 1673] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 1674] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1675] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 1676] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 1677] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 1678] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 1679] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1680] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1681] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 1682] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1683] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 1684] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1685] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1686] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1687] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1688] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 1689] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1690] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1691] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 1692] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 1693] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1694] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1695] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 1696] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1697] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 1698] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1699] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 1700] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 1701] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1702] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 1703] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 1704] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 1705] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1706] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 1707] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 1708] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 1709] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1710] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 1711] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1712] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1713] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 1714] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1715] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 1716] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1717] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 1718] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1719] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 1720] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 1721] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1722] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1723] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 1724] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1725] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 1726] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1727] = 32'b01000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 1728] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1729] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 1730] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 1731] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1732] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[ 1733] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 1734] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1735] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1736] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 1737] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 1738] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1739] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 1740] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 1741] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 1742] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1743] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 1744] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 1745] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1746] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 1747] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 1748] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 1749] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 1750] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 1751] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 1752] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1753] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1754] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1755] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1756] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1757] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 1758] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 1759] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 1760] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 1761] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 1762] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 1763] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 1764] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 1765] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 1766] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1767] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 1768] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 1769] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 1770] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1771] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 1772] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 1773] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1774] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 1775] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 1776] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 1777] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 1778] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 1779] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1780] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 1781] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 1782] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1783] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1784] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1785] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 1786] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 1787] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 1788] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1789] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 1790] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1791] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 1792] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 1793] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1794] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 1795] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1796] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 1797] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 1798] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 1799] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 1800] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 1801] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1802] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 1803] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1804] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 1805] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 1806] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1807] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 1808] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1809] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1810] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 1811] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1812] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1813] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 1814] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 1815] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 1816] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 1817] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 1818] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 1819] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 1820] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 1821] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1822] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 1823] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1824] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1825] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 1826] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 1827] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1828] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1829] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 1830] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1831] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 1832] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 1833] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 1834] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 1835] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1836] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 1837] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1838] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 1839] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1840] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 1841] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 1842] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1843] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1844] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 1845] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1846] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1847] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 1848] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 1849] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1850] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 1851] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 1852] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 1853] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1854] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1855] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 1856] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 1857] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 1858] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1859] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 1860] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1861] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1862] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 1863] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1864] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 1865] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1866] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1867] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 1868] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 1869] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 1870] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1871] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1872] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 1873] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1874] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 1875] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 1876] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 1877] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 1878] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1879] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 1880] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1881] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1882] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1883] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 1884] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 1885] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 1886] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 1887] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 1888] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 1889] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 1890] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 1891] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 1892] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 1893] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1894] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 1895] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 1896] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1897] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 1898] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 1899] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 1900] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1901] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 1902] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 1903] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1904] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 1905] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 1906] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 1907] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 1908] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 1909] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 1910] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 1911] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 1912] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1913] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 1914] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 1915] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 1916] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1917] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1918] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 1919] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1920] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1921] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 1922] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 1923] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1924] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1925] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 1926] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 1927] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1928] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1929] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 1930] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1931] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 1932] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 1933] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 1934] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1935] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 1936] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 1937] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1938] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1939] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 1940] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1941] = 32'b01000010111001100000000000000000;
	assign	noise_gru_input_weights_array[ 1942] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1943] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 1944] = 32'b11000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 1945] = 32'b01000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 1946] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 1947] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1948] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 1949] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 1950] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1951] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1952] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 1953] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 1954] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1955] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 1956] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 1957] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 1958] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 1959] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 1960] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 1961] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 1962] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1963] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 1964] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 1965] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 1966] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 1967] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 1968] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 1969] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 1970] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 1971] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 1972] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 1973] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 1974] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 1975] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1976] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 1977] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 1978] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 1979] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 1980] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 1981] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1982] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 1983] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 1984] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 1985] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 1986] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 1987] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 1988] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 1989] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 1990] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 1991] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 1992] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 1993] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 1994] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1995] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 1996] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 1997] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 1998] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 1999] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2000] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2001] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 2002] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2003] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 2004] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 2005] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2006] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 2007] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2008] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2009] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2010] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2011] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2012] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 2013] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2014] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2015] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 2016] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 2017] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 2018] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2019] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2020] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 2021] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2022] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 2023] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2024] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2025] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 2026] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2027] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2028] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2029] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2030] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 2031] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 2032] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 2033] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2034] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2035] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 2036] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 2037] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2038] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 2039] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2040] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 2041] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2042] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 2043] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 2044] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2045] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2046] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2047] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 2048] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2049] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 2050] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 2051] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2052] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2053] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 2054] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2055] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2056] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 2057] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 2058] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2059] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 2060] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 2061] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2062] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2063] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 2064] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2065] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 2066] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2067] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 2068] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 2069] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 2070] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2071] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 2072] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2073] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2074] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 2075] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2076] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 2077] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 2078] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 2079] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2080] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2081] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2082] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2083] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2084] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2085] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 2086] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2087] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 2088] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 2089] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2090] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 2091] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 2092] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 2093] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 2094] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2095] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 2096] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2097] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2098] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2099] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 2100] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2101] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2102] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2103] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2104] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 2105] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2106] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 2107] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 2108] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 2109] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 2110] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2111] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 2112] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2113] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 2114] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2115] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2116] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 2117] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2118] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 2119] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 2120] = 32'b01000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 2121] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2122] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2123] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 2124] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2125] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 2126] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 2127] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2128] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 2129] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 2130] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 2131] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 2132] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 2133] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 2134] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 2135] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 2136] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 2137] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2138] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 2139] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2140] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 2141] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2142] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 2143] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2144] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2145] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2146] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2147] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2148] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 2149] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 2150] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2151] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2152] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2153] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 2154] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 2155] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 2156] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 2157] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 2158] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2159] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 2160] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 2161] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 2162] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2163] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 2164] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 2165] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 2166] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 2167] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2168] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 2169] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 2170] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 2171] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 2172] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2173] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2174] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 2175] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 2176] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2177] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2178] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 2179] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 2180] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 2181] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 2182] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2183] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2184] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 2185] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 2186] = 32'b11000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 2187] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 2188] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2189] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 2190] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 2191] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 2192] = 32'b01000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 2193] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2194] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2195] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2196] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2197] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 2198] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2199] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2200] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 2201] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 2202] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 2203] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 2204] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 2205] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2206] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 2207] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 2208] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 2209] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 2210] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2211] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2212] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 2213] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 2214] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 2215] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2216] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2217] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2218] = 32'b01000010110111000000000000000000;
	assign	noise_gru_input_weights_array[ 2219] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 2220] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 2221] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2222] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 2223] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2224] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 2225] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 2226] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2227] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 2228] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2229] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2230] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 2231] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 2232] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 2233] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2234] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 2235] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 2236] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 2237] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2238] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 2239] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 2240] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2241] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2242] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 2243] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2244] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2245] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2246] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2247] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 2248] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 2249] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 2250] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2251] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 2252] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 2253] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 2254] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 2255] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2256] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2257] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 2258] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 2259] = 32'b01000010111001100000000000000000;
	assign	noise_gru_input_weights_array[ 2260] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2261] = 32'b11000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 2262] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 2263] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 2264] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 2265] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 2266] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 2267] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 2268] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 2269] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2270] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 2271] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2272] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2273] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2274] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2275] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2276] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2277] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2278] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 2279] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2280] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 2281] = 32'b11000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 2282] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 2283] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2284] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 2285] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 2286] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2287] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 2288] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 2289] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 2290] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 2291] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 2292] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2293] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2294] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 2295] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 2296] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2297] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 2298] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 2299] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2300] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 2301] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 2302] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2303] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 2304] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2305] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2306] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2307] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 2308] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2309] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2310] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2311] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 2312] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 2313] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 2314] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2315] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 2316] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 2317] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2318] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 2319] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2320] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2321] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 2322] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2323] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2324] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 2325] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 2326] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2327] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2328] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2329] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2330] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 2331] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 2332] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2333] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 2334] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2335] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2336] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 2337] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 2338] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 2339] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2340] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2341] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2342] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2343] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2344] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2345] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2346] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2347] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2348] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 2349] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 2350] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2351] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 2352] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 2353] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2354] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 2355] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2356] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 2357] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 2358] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 2359] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 2360] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 2361] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2362] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2363] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2364] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 2365] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 2366] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2367] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2368] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 2369] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 2370] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2371] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 2372] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2373] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 2374] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 2375] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 2376] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 2377] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 2378] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2379] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 2380] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2381] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2382] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 2383] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 2384] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 2385] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 2386] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 2387] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2388] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 2389] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 2390] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 2391] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 2392] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 2393] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 2394] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 2395] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2396] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 2397] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 2398] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 2399] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 2400] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 2401] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 2402] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 2403] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2404] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2405] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2406] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2407] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 2408] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2409] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2410] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 2411] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2412] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2413] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 2414] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2415] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2416] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 2417] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 2418] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 2419] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2420] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2421] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 2422] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 2423] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2424] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 2425] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2426] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2427] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 2428] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2429] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 2430] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 2431] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2432] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 2433] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 2434] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2435] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 2436] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 2437] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 2438] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2439] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 2440] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 2441] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 2442] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 2443] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2444] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 2445] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 2446] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 2447] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 2448] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 2449] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2450] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2451] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2452] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2453] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2454] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2455] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2456] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 2457] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2458] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 2459] = 32'b01000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 2460] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 2461] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2462] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 2463] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 2464] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2465] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 2466] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2467] = 32'b11000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 2468] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2469] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 2470] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2471] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2472] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2473] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 2474] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 2475] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 2476] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2477] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2478] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 2479] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2480] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2481] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 2482] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2483] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 2484] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2485] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 2486] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 2487] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 2488] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 2489] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 2490] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 2491] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2492] = 32'b01000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 2493] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 2494] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 2495] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 2496] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 2497] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 2498] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2499] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 2500] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 2501] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 2502] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 2503] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 2504] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2505] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2506] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 2507] = 32'b11000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 2508] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 2509] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 2510] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2511] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 2512] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2513] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 2514] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2515] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 2516] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 2517] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2518] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 2519] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 2520] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 2521] = 32'b11000010110010100000000000000000;
	assign	noise_gru_input_weights_array[ 2522] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 2523] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2524] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2525] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2526] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 2527] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 2528] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 2529] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 2530] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 2531] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 2532] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 2533] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2534] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 2535] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2536] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2537] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 2538] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 2539] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 2540] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 2541] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 2542] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 2543] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2544] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 2545] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2546] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2547] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 2548] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2549] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2550] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 2551] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2552] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 2553] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 2554] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 2555] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2556] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2557] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2558] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 2559] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2560] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 2561] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 2562] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2563] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 2564] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2565] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 2566] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 2567] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 2568] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2569] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 2570] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 2571] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2572] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 2573] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 2574] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 2575] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 2576] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2577] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 2578] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 2579] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 2580] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2581] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2582] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2583] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 2584] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2585] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 2586] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 2587] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 2588] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 2589] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 2590] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2591] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 2592] = 32'b01000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2593] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 2594] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2595] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2596] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 2597] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 2598] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2599] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2600] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 2601] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 2602] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 2603] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 2604] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2605] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 2606] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 2607] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2608] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 2609] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 2610] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 2611] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2612] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2613] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2614] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2615] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 2616] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2617] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 2618] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 2619] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2620] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2621] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2622] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 2623] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2624] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 2625] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2626] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2627] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2628] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 2629] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2630] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 2631] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 2632] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2633] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 2634] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 2635] = 32'b01000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 2636] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2637] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2638] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2639] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 2640] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 2641] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 2642] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 2643] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2644] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 2645] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2646] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 2647] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 2648] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 2649] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2650] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 2651] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 2652] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2653] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 2654] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 2655] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 2656] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2657] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 2658] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 2659] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 2660] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 2661] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 2662] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2663] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2664] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2665] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 2666] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2667] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 2668] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2669] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2670] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[ 2671] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2672] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 2673] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2674] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 2675] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 2676] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 2677] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 2678] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 2679] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2680] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 2681] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 2682] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2683] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2684] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 2685] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 2686] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 2687] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 2688] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 2689] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2690] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 2691] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 2692] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 2693] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 2694] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 2695] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2696] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 2697] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 2698] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2699] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2700] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2701] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 2702] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 2703] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2704] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 2705] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 2706] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2707] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2708] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 2709] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 2710] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2711] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2712] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 2713] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2714] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 2715] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 2716] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 2717] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 2718] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2719] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 2720] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 2721] = 32'b01000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 2722] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2723] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 2724] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2725] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2726] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 2727] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2728] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2729] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 2730] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2731] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2732] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2733] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 2734] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2735] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2736] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2737] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2738] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 2739] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 2740] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 2741] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2742] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 2743] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2744] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2745] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2746] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2747] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 2748] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 2749] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2750] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2751] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 2752] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2753] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 2754] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2755] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 2756] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 2757] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 2758] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 2759] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2760] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2761] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 2762] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2763] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2764] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 2765] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 2766] = 32'b01000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 2767] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 2768] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[ 2769] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 2770] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2771] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 2772] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2773] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2774] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 2775] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 2776] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[ 2777] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2778] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 2779] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2780] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 2781] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 2782] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 2783] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 2784] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 2785] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 2786] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2787] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2788] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2789] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 2790] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 2791] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2792] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2793] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 2794] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 2795] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 2796] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 2797] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 2798] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 2799] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 2800] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2801] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 2802] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2803] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2804] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 2805] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 2806] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2807] = 32'b01000010111001100000000000000000;
	assign	noise_gru_input_weights_array[ 2808] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 2809] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 2810] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 2811] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2812] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 2813] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 2814] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2815] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 2816] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 2817] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2818] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 2819] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2820] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 2821] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 2822] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 2823] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2824] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2825] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 2826] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2827] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2828] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 2829] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 2830] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2831] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 2832] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 2833] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 2834] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 2835] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2836] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 2837] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 2838] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 2839] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 2840] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2841] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 2842] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2843] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 2844] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2845] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2846] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2847] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 2848] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 2849] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 2850] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 2851] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 2852] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 2853] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 2854] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 2855] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 2856] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2857] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 2858] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 2859] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 2860] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2861] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 2862] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2863] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2864] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2865] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 2866] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 2867] = 32'b01000010110111000000000000000000;
	assign	noise_gru_input_weights_array[ 2868] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2869] = 32'b01000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 2870] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2871] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 2872] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2873] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 2874] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 2875] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2876] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 2877] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 2878] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 2879] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 2880] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 2881] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2882] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2883] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 2884] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 2885] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2886] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 2887] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 2888] = 32'b11000010110111000000000000000000;
	assign	noise_gru_input_weights_array[ 2889] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 2890] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2891] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 2892] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 2893] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2894] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 2895] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 2896] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 2897] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 2898] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 2899] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 2900] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2901] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 2902] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2903] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 2904] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2905] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 2906] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 2907] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 2908] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 2909] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2910] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2911] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 2912] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2913] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2914] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2915] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 2916] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 2917] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 2918] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2919] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2920] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2921] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2922] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2923] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 2924] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 2925] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 2926] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2927] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 2928] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2929] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2930] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2931] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2932] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2933] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2934] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 2935] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[ 2936] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2937] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2938] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2939] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2940] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2941] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2942] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 2943] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 2944] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 2945] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 2946] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2947] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2948] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 2949] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 2950] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 2951] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 2952] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 2953] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 2954] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 2955] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2956] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2957] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 2958] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 2959] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 2960] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 2961] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 2962] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 2963] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 2964] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2965] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 2966] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 2967] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 2968] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 2969] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 2970] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 2971] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2972] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 2973] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 2974] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 2975] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 2976] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 2977] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 2978] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 2979] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 2980] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 2981] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 2982] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 2983] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 2984] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2985] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 2986] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 2987] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 2988] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 2989] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 2990] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 2991] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 2992] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 2993] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 2994] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 2995] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 2996] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 2997] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 2998] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 2999] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 3000] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 3001] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3002] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 3003] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 3004] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 3005] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3006] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3007] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 3008] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 3009] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3010] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3011] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 3012] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3013] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3014] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3015] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 3016] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 3017] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 3018] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 3019] = 32'b11000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 3020] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 3021] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 3022] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 3023] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 3024] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 3025] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 3026] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3027] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 3028] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3029] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3030] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3031] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3032] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3033] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3034] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 3035] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 3036] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 3037] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3038] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 3039] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3040] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3041] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 3042] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 3043] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 3044] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 3045] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 3046] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3047] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 3048] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 3049] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 3050] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3051] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3052] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 3053] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3054] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3055] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3056] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 3057] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3058] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3059] = 32'b11000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 3060] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3061] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 3062] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 3063] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 3064] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 3065] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 3066] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 3067] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 3068] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3069] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 3070] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3071] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 3072] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 3073] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3074] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3075] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 3076] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 3077] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 3078] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 3079] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 3080] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3081] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3082] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3083] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 3084] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3085] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 3086] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3087] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 3088] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3089] = 32'b01000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 3090] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3091] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3092] = 32'b11000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 3093] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3094] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 3095] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 3096] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 3097] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 3098] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 3099] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3100] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 3101] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 3102] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3103] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 3104] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 3105] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 3106] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 3107] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 3108] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3109] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 3110] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3111] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3112] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3113] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3114] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 3115] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3116] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3117] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 3118] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 3119] = 32'b11000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 3120] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 3121] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 3122] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 3123] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3124] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 3125] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 3126] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 3127] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 3128] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 3129] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3130] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3131] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 3132] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 3133] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3134] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 3135] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3136] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 3137] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 3138] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 3139] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3140] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3141] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 3142] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 3143] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 3144] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3145] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3146] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3147] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3148] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 3149] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 3150] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 3151] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3152] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 3153] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3154] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3155] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 3156] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 3157] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 3158] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 3159] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3160] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 3161] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 3162] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 3163] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 3164] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3165] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 3166] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 3167] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 3168] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 3169] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 3170] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3171] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 3172] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3173] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 3174] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 3175] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3176] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 3177] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 3178] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3179] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3180] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3181] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 3182] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3183] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 3184] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 3185] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3186] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3187] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 3188] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 3189] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3190] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3191] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3192] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 3193] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3194] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 3195] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3196] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3197] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3198] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 3199] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 3200] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 3201] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 3202] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3203] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 3204] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 3205] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 3206] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3207] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 3208] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 3209] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3210] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 3211] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 3212] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 3213] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3214] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 3215] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 3216] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 3217] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 3218] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 3219] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 3220] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 3221] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3222] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3223] = 32'b11000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 3224] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 3225] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 3226] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 3227] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 3228] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 3229] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3230] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 3231] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 3232] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3233] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 3234] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 3235] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 3236] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3237] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3238] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3239] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3240] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 3241] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 3242] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3243] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3244] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 3245] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 3246] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 3247] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 3248] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3249] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 3250] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 3251] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 3252] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 3253] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3254] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 3255] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 3256] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3257] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 3258] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 3259] = 32'b11000010110010100000000000000000;
	assign	noise_gru_input_weights_array[ 3260] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 3261] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 3262] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 3263] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 3264] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3265] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 3266] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 3267] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 3268] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 3269] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 3270] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 3271] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 3272] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3273] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 3274] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3275] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3276] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3277] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 3278] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 3279] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 3280] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3281] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 3282] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 3283] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 3284] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 3285] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3286] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3287] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 3288] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3289] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 3290] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 3291] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3292] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 3293] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3294] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3295] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 3296] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 3297] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 3298] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3299] = 32'b01000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 3300] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 3301] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 3302] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3303] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 3304] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3305] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3306] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3307] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 3308] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3309] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 3310] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 3311] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3312] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 3313] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3314] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 3315] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 3316] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3317] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3318] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 3319] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3320] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 3321] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3322] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 3323] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 3324] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3325] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3326] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3327] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 3328] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3329] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3330] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 3331] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3332] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 3333] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3334] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 3335] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 3336] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 3337] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 3338] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 3339] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 3340] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 3341] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 3342] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3343] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3344] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 3345] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3346] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 3347] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 3348] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3349] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3350] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3351] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3352] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3353] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 3354] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 3355] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3356] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 3357] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 3358] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 3359] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 3360] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3361] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 3362] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 3363] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3364] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 3365] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 3366] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3367] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 3368] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 3369] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3370] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 3371] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3372] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 3373] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 3374] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 3375] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 3376] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3377] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3378] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3379] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 3380] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 3381] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 3382] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3383] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 3384] = 32'b11000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 3385] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3386] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 3387] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 3388] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3389] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 3390] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3391] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 3392] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3393] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3394] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 3395] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 3396] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3397] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 3398] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3399] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 3400] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3401] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3402] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 3403] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 3404] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 3405] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 3406] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 3407] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 3408] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3409] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3410] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 3411] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3412] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3413] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 3414] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 3415] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3416] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 3417] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 3418] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3419] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 3420] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3421] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3422] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 3423] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 3424] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 3425] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3426] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3427] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3428] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3429] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 3430] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 3431] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 3432] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 3433] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 3434] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 3435] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 3436] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 3437] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 3438] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 3439] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 3440] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 3441] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 3442] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 3443] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3444] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 3445] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 3446] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 3447] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 3448] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 3449] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 3450] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 3451] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3452] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3453] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3454] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 3455] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 3456] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 3457] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3458] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3459] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 3460] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3461] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3462] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 3463] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 3464] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 3465] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3466] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3467] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 3468] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3469] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 3470] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 3471] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 3472] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3473] = 32'b01000010111001100000000000000000;
	assign	noise_gru_input_weights_array[ 3474] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 3475] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 3476] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 3477] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 3478] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 3479] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 3480] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3481] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3482] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3483] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 3484] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3485] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3486] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3487] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 3488] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 3489] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 3490] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3491] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3492] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 3493] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 3494] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 3495] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3496] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 3497] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 3498] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 3499] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 3500] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3501] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 3502] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 3503] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 3504] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 3505] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3506] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 3507] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3508] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3509] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3510] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3511] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 3512] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 3513] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3514] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3515] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 3516] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 3517] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 3518] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 3519] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3520] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3521] = 32'b11000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 3522] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 3523] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 3524] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3525] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 3526] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 3527] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3528] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 3529] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3530] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 3531] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 3532] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 3533] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 3534] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 3535] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3536] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 3537] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3538] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 3539] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 3540] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3541] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 3542] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3543] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3544] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3545] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 3546] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3547] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3548] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 3549] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 3550] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 3551] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3552] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 3553] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3554] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 3555] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3556] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3557] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 3558] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 3559] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 3560] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 3561] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3562] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3563] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 3564] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 3565] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3566] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3567] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 3568] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 3569] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 3570] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3571] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 3572] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 3573] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 3574] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 3575] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3576] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 3577] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3578] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3579] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 3580] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3581] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3582] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3583] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 3584] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3585] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3586] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3587] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 3588] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 3589] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 3590] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 3591] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 3592] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 3593] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3594] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 3595] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3596] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3597] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3598] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 3599] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3600] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 3601] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 3602] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 3603] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 3604] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3605] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3606] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3607] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 3608] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 3609] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 3610] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3611] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3612] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3613] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3614] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 3615] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 3616] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 3617] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 3618] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3619] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 3620] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 3621] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 3622] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3623] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3624] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 3625] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3626] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3627] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3628] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 3629] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 3630] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 3631] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 3632] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 3633] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 3634] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3635] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 3636] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3637] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 3638] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 3639] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3640] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3641] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3642] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 3643] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 3644] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 3645] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 3646] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3647] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 3648] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 3649] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 3650] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3651] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3652] = 32'b11000010110111000000000000000000;
	assign	noise_gru_input_weights_array[ 3653] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 3654] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 3655] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 3656] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 3657] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 3658] = 32'b11000010110111000000000000000000;
	assign	noise_gru_input_weights_array[ 3659] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 3660] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3661] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3662] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3663] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 3664] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 3665] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 3666] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3667] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 3668] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3669] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3670] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3671] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 3672] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 3673] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3674] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3675] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3676] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 3677] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 3678] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 3679] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 3680] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3681] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3682] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3683] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 3684] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 3685] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 3686] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3687] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 3688] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 3689] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 3690] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3691] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 3692] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 3693] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3694] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 3695] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3696] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3697] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 3698] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 3699] = 32'b11000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 3700] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3701] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 3702] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3703] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 3704] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 3705] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 3706] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 3707] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 3708] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3709] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 3710] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 3711] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 3712] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 3713] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3714] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3715] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 3716] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3717] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3718] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3719] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3720] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 3721] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 3722] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3723] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3724] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3725] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 3726] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3727] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3728] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3729] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 3730] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 3731] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 3732] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 3733] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 3734] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3735] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3736] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 3737] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 3738] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3739] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 3740] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3741] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3742] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 3743] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 3744] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 3745] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 3746] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 3747] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3748] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 3749] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3750] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3751] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 3752] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 3753] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 3754] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 3755] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 3756] = 32'b11000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 3757] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 3758] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 3759] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3760] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3761] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3762] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3763] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 3764] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 3765] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 3766] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 3767] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3768] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3769] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3770] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3771] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3772] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 3773] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 3774] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3775] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 3776] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3777] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3778] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 3779] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3780] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 3781] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3782] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 3783] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 3784] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 3785] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 3786] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 3787] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 3788] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 3789] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 3790] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 3791] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 3792] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 3793] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 3794] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 3795] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3796] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 3797] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 3798] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3799] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3800] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3801] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 3802] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 3803] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3804] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 3805] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 3806] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3807] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3808] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 3809] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 3810] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3811] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 3812] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 3813] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 3814] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 3815] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 3816] = 32'b11000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 3817] = 32'b01000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3818] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3819] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 3820] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 3821] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3822] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 3823] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 3824] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 3825] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 3826] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 3827] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 3828] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 3829] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3830] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 3831] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 3832] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 3833] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 3834] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 3835] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3836] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3837] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 3838] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 3839] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 3840] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3841] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 3842] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3843] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3844] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3845] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3846] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3847] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 3848] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 3849] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 3850] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 3851] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 3852] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 3853] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 3854] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3855] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 3856] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 3857] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3858] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3859] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 3860] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 3861] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3862] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 3863] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3864] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 3865] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 3866] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 3867] = 32'b11000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 3868] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3869] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 3870] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 3871] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 3872] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3873] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3874] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 3875] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3876] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 3877] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3878] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 3879] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3880] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3881] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 3882] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3883] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3884] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3885] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 3886] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 3887] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3888] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 3889] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 3890] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3891] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3892] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 3893] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 3894] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3895] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 3896] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 3897] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3898] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 3899] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 3900] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3901] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 3902] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3903] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 3904] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 3905] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 3906] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3907] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3908] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 3909] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 3910] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 3911] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3912] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 3913] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3914] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3915] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 3916] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3917] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 3918] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 3919] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3920] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3921] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3922] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3923] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 3924] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 3925] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 3926] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 3927] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 3928] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 3929] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 3930] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3931] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3932] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3933] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 3934] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3935] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 3936] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 3937] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 3938] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 3939] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 3940] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3941] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 3942] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 3943] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3944] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 3945] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 3946] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 3947] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 3948] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 3949] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3950] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 3951] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 3952] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 3953] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3954] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3955] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 3956] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3957] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3958] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 3959] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 3960] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 3961] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3962] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 3963] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 3964] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 3965] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 3966] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 3967] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3968] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3969] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 3970] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 3971] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 3972] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 3973] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 3974] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3975] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 3976] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 3977] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 3978] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 3979] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 3980] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 3981] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 3982] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 3983] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 3984] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3985] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 3986] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 3987] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3988] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 3989] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 3990] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 3991] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 3992] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 3993] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 3994] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 3995] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 3996] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 3997] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 3998] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 3999] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 4000] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 4001] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4002] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 4003] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 4004] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 4005] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 4006] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 4007] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4008] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4009] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 4010] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4011] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 4012] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4013] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4014] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 4015] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 4016] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4017] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 4018] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 4019] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4020] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4021] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 4022] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 4023] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 4024] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 4025] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4026] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4027] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 4028] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4029] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4030] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 4031] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4032] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 4033] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4034] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 4035] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 4036] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4037] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4038] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 4039] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 4040] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 4041] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4042] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4043] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 4044] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 4045] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4046] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4047] = 32'b01000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 4048] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 4049] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4050] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 4051] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 4052] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 4053] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 4054] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4055] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4056] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 4057] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4058] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4059] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4060] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4061] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4062] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 4063] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 4064] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4065] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 4066] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4067] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 4068] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4069] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4070] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 4071] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 4072] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4073] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4074] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 4075] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4076] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 4077] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4078] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 4079] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4080] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4081] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4082] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 4083] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 4084] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4085] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 4086] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4087] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4088] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4089] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 4090] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 4091] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 4092] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 4093] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 4094] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 4095] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4096] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 4097] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 4098] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 4099] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 4100] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 4101] = 32'b11000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 4102] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 4103] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 4104] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 4105] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4106] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 4107] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4108] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4109] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 4110] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 4111] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4112] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4113] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 4114] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 4115] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 4116] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 4117] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[ 4118] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 4119] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 4120] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 4121] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 4122] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 4123] = 32'b11000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 4124] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 4125] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 4126] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4127] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4128] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 4129] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4130] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4131] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 4132] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 4133] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 4134] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4135] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4136] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4137] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 4138] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4139] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 4140] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 4141] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4142] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4143] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 4144] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4145] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4146] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 4147] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4148] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 4149] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 4150] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 4151] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4152] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 4153] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 4154] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4155] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 4156] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4157] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 4158] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4159] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4160] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4161] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 4162] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4163] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4164] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4165] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 4166] = 32'b11000010110010100000000000000000;
	assign	noise_gru_input_weights_array[ 4167] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[ 4168] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4169] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4170] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4171] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 4172] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 4173] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4174] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 4175] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 4176] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 4177] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 4178] = 32'b01000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 4179] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 4180] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4181] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4182] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4183] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 4184] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 4185] = 32'b01000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4186] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4187] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4188] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 4189] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 4190] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4191] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 4192] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 4193] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4194] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 4195] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 4196] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4197] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4198] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4199] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 4200] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4201] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 4202] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4203] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 4204] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4205] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4206] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4207] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 4208] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 4209] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 4210] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4211] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 4212] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 4213] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 4214] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 4215] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 4216] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 4217] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4218] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4219] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 4220] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 4221] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4222] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4223] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4224] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 4225] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 4226] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4227] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 4228] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 4229] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 4230] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4231] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4232] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4233] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4234] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 4235] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 4236] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 4237] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 4238] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4239] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4240] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 4241] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4242] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4243] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4244] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 4245] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 4246] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4247] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 4248] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4249] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4250] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4251] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4252] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4253] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4254] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 4255] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 4256] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4257] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 4258] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 4259] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4260] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4261] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4262] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4263] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 4264] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 4265] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 4266] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 4267] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4268] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4269] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 4270] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4271] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 4272] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4273] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4274] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4275] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 4276] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4277] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 4278] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 4279] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 4280] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4281] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4282] = 32'b01000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 4283] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 4284] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 4285] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4286] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 4287] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4288] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 4289] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 4290] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 4291] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 4292] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4293] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4294] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4295] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 4296] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4297] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4298] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 4299] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 4300] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 4301] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 4302] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 4303] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 4304] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 4305] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 4306] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 4307] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 4308] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4309] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4310] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 4311] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 4312] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 4313] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4314] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4315] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4316] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4317] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4318] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 4319] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 4320] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 4321] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4322] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4323] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 4324] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 4325] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4326] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4327] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 4328] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 4329] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4330] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 4331] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 4332] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4333] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4334] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4335] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 4336] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4337] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4338] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 4339] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 4340] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4341] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4342] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 4343] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 4344] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 4345] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4346] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4347] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4348] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4349] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 4350] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4351] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4352] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 4353] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 4354] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4355] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4356] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4357] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4358] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4359] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 4360] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 4361] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4362] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 4363] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4364] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4365] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 4366] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4367] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 4368] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4369] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 4370] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 4371] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4372] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4373] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 4374] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4375] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4376] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 4377] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 4378] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 4379] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4380] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 4381] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 4382] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 4383] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 4384] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 4385] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 4386] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 4387] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 4388] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 4389] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 4390] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 4391] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4392] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4393] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 4394] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 4395] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 4396] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4397] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 4398] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 4399] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 4400] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 4401] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4402] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 4403] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 4404] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 4405] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 4406] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 4407] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 4408] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 4409] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 4410] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 4411] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4412] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4413] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4414] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 4415] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 4416] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 4417] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4418] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 4419] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 4420] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 4421] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 4422] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 4423] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 4424] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 4425] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 4426] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 4427] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 4428] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4429] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 4430] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4431] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 4432] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 4433] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4434] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 4435] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4436] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 4437] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 4438] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 4439] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4440] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4441] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 4442] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 4443] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 4444] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 4445] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 4446] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4447] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 4448] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 4449] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4450] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4451] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 4452] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 4453] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4454] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 4455] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4456] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4457] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 4458] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4459] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4460] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4461] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 4462] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 4463] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4464] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 4465] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 4466] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4467] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 4468] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 4469] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4470] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 4471] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4472] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 4473] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4474] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 4475] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 4476] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4477] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 4478] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 4479] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4480] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4481] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 4482] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4483] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4484] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 4485] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 4486] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4487] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 4488] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 4489] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 4490] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 4491] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 4492] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 4493] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4494] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 4495] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 4496] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4497] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 4498] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4499] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4500] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 4501] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4502] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4503] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4504] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 4505] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4506] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 4507] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4508] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4509] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4510] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4511] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 4512] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 4513] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4514] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 4515] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4516] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 4517] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4518] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4519] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 4520] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 4521] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4522] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 4523] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4524] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4525] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 4526] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 4527] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4528] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 4529] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 4530] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4531] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 4532] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4533] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 4534] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4535] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 4536] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4537] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 4538] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4539] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 4540] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 4541] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 4542] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4543] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 4544] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 4545] = 32'b01000010110111000000000000000000;
	assign	noise_gru_input_weights_array[ 4546] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4547] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 4548] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 4549] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 4550] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4551] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4552] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4553] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4554] = 32'b11000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 4555] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 4556] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 4557] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 4558] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 4559] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 4560] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4561] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 4562] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4563] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4564] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4565] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4566] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4567] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 4568] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 4569] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 4570] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 4571] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4572] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4573] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4574] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 4575] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 4576] = 32'b01000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4577] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 4578] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4579] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4580] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4581] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 4582] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4583] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4584] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4585] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 4586] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 4587] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 4588] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 4589] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 4590] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 4591] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 4592] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 4593] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 4594] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 4595] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 4596] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 4597] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 4598] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4599] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 4600] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4601] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 4602] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 4603] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 4604] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 4605] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 4606] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 4607] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 4608] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4609] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4610] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4611] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4612] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4613] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 4614] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 4615] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 4616] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 4617] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4618] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 4619] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 4620] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 4621] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 4622] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 4623] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4624] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 4625] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 4626] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4627] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4628] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 4629] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4630] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 4631] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 4632] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4633] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4634] = 32'b11000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 4635] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 4636] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4637] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 4638] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 4639] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 4640] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4641] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4642] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 4643] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 4644] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4645] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4646] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 4647] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4648] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4649] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4650] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 4651] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 4652] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4653] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 4654] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4655] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 4656] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 4657] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4658] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4659] = 32'b11000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 4660] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 4661] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 4662] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4663] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4664] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4665] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4666] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 4667] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4668] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4669] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4670] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4671] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[ 4672] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4673] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4674] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4675] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 4676] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 4677] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4678] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 4679] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4680] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 4681] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 4682] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 4683] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 4684] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4685] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 4686] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4687] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 4688] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4689] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 4690] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 4691] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 4692] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 4693] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4694] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4695] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4696] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4697] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4698] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 4699] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4700] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4701] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 4702] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 4703] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 4704] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4705] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 4706] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4707] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 4708] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4709] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4710] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4711] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4712] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4713] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4714] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 4715] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 4716] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4717] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4718] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4719] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4720] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4721] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 4722] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4723] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4724] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 4725] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 4726] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4727] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 4728] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4729] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4730] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 4731] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4732] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 4733] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4734] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4735] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4736] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 4737] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 4738] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 4739] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 4740] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4741] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4742] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4743] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 4744] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4745] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 4746] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4747] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 4748] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 4749] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4750] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4751] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4752] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 4753] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4754] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4755] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 4756] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4757] = 32'b01000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 4758] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 4759] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[ 4760] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 4761] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 4762] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 4763] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 4764] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 4765] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4766] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4767] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 4768] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4769] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 4770] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 4771] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4772] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 4773] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4774] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 4775] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4776] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4777] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4778] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4779] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4780] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4781] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4782] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 4783] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4784] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 4785] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 4786] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 4787] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 4788] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 4789] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 4790] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 4791] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 4792] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 4793] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 4794] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 4795] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4796] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4797] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4798] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 4799] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 4800] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4801] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 4802] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4803] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 4804] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4805] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 4806] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4807] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 4808] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 4809] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 4810] = 32'b11000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 4811] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 4812] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4813] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 4814] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4815] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 4816] = 32'b01000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4817] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4818] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 4819] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4820] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 4821] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 4822] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4823] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4824] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 4825] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 4826] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4827] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 4828] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4829] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4830] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 4831] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4832] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 4833] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4834] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 4835] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 4836] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 4837] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4838] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 4839] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 4840] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 4841] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 4842] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 4843] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 4844] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4845] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 4846] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 4847] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4848] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4849] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4850] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4851] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 4852] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4853] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4854] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4855] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 4856] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4857] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 4858] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 4859] = 32'b11000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 4860] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 4861] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 4862] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4863] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4864] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 4865] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 4866] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4867] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 4868] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4869] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4870] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4871] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4872] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4873] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 4874] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 4875] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 4876] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4877] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 4878] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 4879] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 4880] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4881] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 4882] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4883] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 4884] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 4885] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4886] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 4887] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 4888] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4889] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4890] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4891] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4892] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 4893] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4894] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 4895] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4896] = 32'b11000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 4897] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4898] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 4899] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 4900] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4901] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4902] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4903] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4904] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 4905] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 4906] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4907] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 4908] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4909] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4910] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4911] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4912] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 4913] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4914] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 4915] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 4916] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4917] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 4918] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 4919] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 4920] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 4921] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 4922] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 4923] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 4924] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 4925] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4926] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4927] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4928] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4929] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 4930] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 4931] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4932] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4933] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 4934] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 4935] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 4936] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 4937] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4938] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 4939] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4940] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 4941] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 4942] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4943] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 4944] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 4945] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4946] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 4947] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4948] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4949] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 4950] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 4951] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 4952] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 4953] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 4954] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 4955] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 4956] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 4957] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 4958] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 4959] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 4960] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 4961] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4962] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4963] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4964] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 4965] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4966] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 4967] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 4968] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 4969] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4970] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4971] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 4972] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 4973] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4974] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 4975] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4976] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 4977] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4978] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4979] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 4980] = 32'b11000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 4981] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4982] = 32'b11000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 4983] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 4984] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 4985] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4986] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 4987] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4988] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4989] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 4990] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 4991] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 4992] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 4993] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 4994] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 4995] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 4996] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4997] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 4998] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 4999] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5000] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 5001] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 5002] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 5003] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5004] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 5005] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5006] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5007] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 5008] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 5009] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5010] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 5011] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5012] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5013] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 5014] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5015] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 5016] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5017] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5018] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5019] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 5020] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 5021] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 5022] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 5023] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5024] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 5025] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5026] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5027] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 5028] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 5029] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 5030] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 5031] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 5032] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 5033] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 5034] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 5035] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5036] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 5037] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 5038] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 5039] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 5040] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5041] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5042] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 5043] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5044] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5045] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 5046] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5047] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 5048] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 5049] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5050] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 5051] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 5052] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5053] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 5054] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 5055] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 5056] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5057] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 5058] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 5059] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5060] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5061] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5062] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5063] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 5064] = 32'b01000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 5065] = 32'b11000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 5066] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5067] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 5068] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 5069] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 5070] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 5071] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5072] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 5073] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5074] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5075] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 5076] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 5077] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 5078] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 5079] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 5080] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 5081] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 5082] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5083] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5084] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 5085] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 5086] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 5087] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 5088] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5089] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 5090] = 32'b01000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5091] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 5092] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 5093] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 5094] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5095] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5096] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5097] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 5098] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 5099] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 5100] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 5101] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 5102] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 5103] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 5104] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 5105] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 5106] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5107] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 5108] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 5109] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 5110] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 5111] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5112] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 5113] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 5114] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5115] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 5116] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 5117] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 5118] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 5119] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5120] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 5121] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5122] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5123] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 5124] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5125] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5126] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 5127] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 5128] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 5129] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5130] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5131] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5132] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 5133] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 5134] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 5135] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 5136] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5137] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5138] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 5139] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 5140] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 5141] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 5142] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5143] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 5144] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 5145] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 5146] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5147] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 5148] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5149] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 5150] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 5151] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 5152] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 5153] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 5154] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 5155] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 5156] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 5157] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5158] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5159] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 5160] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 5161] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 5162] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 5163] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 5164] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 5165] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5166] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 5167] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 5168] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5169] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 5170] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 5171] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5172] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 5173] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 5174] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 5175] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5176] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 5177] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 5178] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5179] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 5180] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 5181] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 5182] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 5183] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 5184] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5185] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 5186] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 5187] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 5188] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 5189] = 32'b01000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5190] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5191] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 5192] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 5193] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5194] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5195] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 5196] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 5197] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 5198] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 5199] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 5200] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 5201] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 5202] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 5203] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 5204] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5205] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 5206] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 5207] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5208] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 5209] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 5210] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 5211] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5212] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 5213] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 5214] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 5215] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 5216] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 5217] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 5218] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5219] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 5220] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5221] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 5222] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5223] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 5224] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 5225] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 5226] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5227] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 5228] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5229] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 5230] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5231] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 5232] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 5233] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 5234] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5235] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 5236] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 5237] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 5238] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5239] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5240] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 5241] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5242] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 5243] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5244] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 5245] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5246] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 5247] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5248] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 5249] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 5250] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 5251] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 5252] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 5253] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5254] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5255] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5256] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 5257] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5258] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 5259] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 5260] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 5261] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 5262] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 5263] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 5264] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5265] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 5266] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 5267] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 5268] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 5269] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5270] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 5271] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 5272] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 5273] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5274] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 5275] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5276] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 5277] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 5278] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5279] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 5280] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 5281] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 5282] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 5283] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 5284] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 5285] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5286] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5287] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5288] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 5289] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 5290] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 5291] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 5292] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 5293] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 5294] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 5295] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 5296] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 5297] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5298] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5299] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5300] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 5301] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5302] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 5303] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 5304] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5305] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 5306] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5307] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 5308] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5309] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 5310] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 5311] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 5312] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5313] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 5314] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 5315] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 5316] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5317] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5318] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5319] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 5320] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5321] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 5322] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 5323] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5324] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5325] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5326] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 5327] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 5328] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 5329] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5330] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 5331] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 5332] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 5333] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 5334] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 5335] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 5336] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 5337] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5338] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 5339] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 5340] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 5341] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 5342] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 5343] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 5344] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 5345] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 5346] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 5347] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 5348] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5349] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 5350] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 5351] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5352] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 5353] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5354] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5355] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5356] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 5357] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 5358] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5359] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 5360] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5361] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 5362] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 5363] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5364] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5365] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 5366] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5367] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5368] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 5369] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5370] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5371] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5372] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 5373] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 5374] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 5375] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 5376] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5377] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 5378] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 5379] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 5380] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 5381] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 5382] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 5383] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 5384] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5385] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 5386] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5387] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 5388] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5389] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5390] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 5391] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 5392] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 5393] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 5394] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 5395] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5396] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 5397] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 5398] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 5399] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 5400] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5401] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 5402] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 5403] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 5404] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 5405] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5406] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5407] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 5408] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 5409] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 5410] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5411] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 5412] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5413] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 5414] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 5415] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 5416] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5417] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 5418] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 5419] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 5420] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 5421] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 5422] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5423] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 5424] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5425] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 5426] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 5427] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5428] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5429] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5430] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5431] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 5432] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 5433] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5434] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 5435] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 5436] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 5437] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 5438] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5439] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5440] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5441] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 5442] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 5443] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 5444] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5445] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 5446] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 5447] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5448] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5449] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5450] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5451] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5452] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 5453] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5454] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5455] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5456] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5457] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5458] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 5459] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 5460] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 5461] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5462] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5463] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 5464] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5465] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 5466] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 5467] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5468] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 5469] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5470] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 5471] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5472] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 5473] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5474] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5475] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 5476] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5477] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 5478] = 32'b11000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 5479] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5480] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 5481] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 5482] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 5483] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5484] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5485] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 5486] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5487] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 5488] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 5489] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5490] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5491] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 5492] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 5493] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5494] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 5495] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5496] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5497] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5498] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5499] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5500] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5501] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5502] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 5503] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 5504] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 5505] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 5506] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 5507] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5508] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5509] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5510] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 5511] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 5512] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 5513] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 5514] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 5515] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 5516] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5517] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5518] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5519] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5520] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 5521] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 5522] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 5523] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 5524] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 5525] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5526] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5527] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 5528] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5529] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5530] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5531] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 5532] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 5533] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 5534] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5535] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 5536] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 5537] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5538] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5539] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 5540] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5541] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 5542] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 5543] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 5544] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5545] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 5546] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 5547] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 5548] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 5549] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5550] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 5551] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5552] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 5553] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5554] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5555] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5556] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5557] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 5558] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5559] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5560] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5561] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5562] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 5563] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5564] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5565] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5566] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 5567] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 5568] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5569] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 5570] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5571] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 5572] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5573] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5574] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5575] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 5576] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5577] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5578] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5579] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 5580] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5581] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5582] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5583] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 5584] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5585] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5586] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5587] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 5588] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 5589] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5590] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 5591] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 5592] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5593] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 5594] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 5595] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 5596] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5597] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5598] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 5599] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 5600] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 5601] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 5602] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 5603] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 5604] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5605] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 5606] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 5607] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5608] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5609] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 5610] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 5611] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5612] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5613] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 5614] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 5615] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5616] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5617] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 5618] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 5619] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 5620] = 32'b11000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 5621] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 5622] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 5623] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 5624] = 32'b11000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 5625] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 5626] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5627] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 5628] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 5629] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 5630] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 5631] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5632] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5633] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5634] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 5635] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 5636] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 5637] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5638] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5639] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5640] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5641] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 5642] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5643] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 5644] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 5645] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 5646] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5647] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5648] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5649] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5650] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 5651] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 5652] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 5653] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 5654] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 5655] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 5656] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 5657] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 5658] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5659] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5660] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 5661] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 5662] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 5663] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 5664] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5665] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5666] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 5667] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5668] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 5669] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 5670] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 5671] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 5672] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5673] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 5674] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 5675] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 5676] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 5677] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 5678] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 5679] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 5680] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 5681] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 5682] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5683] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5684] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 5685] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 5686] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 5687] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 5688] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 5689] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 5690] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 5691] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5692] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5693] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 5694] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 5695] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 5696] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 5697] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 5698] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 5699] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 5700] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5701] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 5702] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 5703] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 5704] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 5705] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5706] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 5707] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 5708] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5709] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 5710] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 5711] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5712] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5713] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5714] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5715] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5716] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5717] = 32'b01000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 5718] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 5719] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5720] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5721] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 5722] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 5723] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5724] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5725] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 5726] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5727] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 5728] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 5729] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 5730] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5731] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 5732] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5733] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 5734] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5735] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5736] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5737] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5738] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 5739] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 5740] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 5741] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 5742] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5743] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 5744] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 5745] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 5746] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 5747] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 5748] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 5749] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 5750] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 5751] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 5752] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 5753] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 5754] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 5755] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 5756] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 5757] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5758] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5759] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 5760] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 5761] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 5762] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 5763] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 5764] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 5765] = 32'b01000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5766] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 5767] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 5768] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 5769] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5770] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 5771] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 5772] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 5773] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 5774] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 5775] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 5776] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 5777] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5778] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5779] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5780] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5781] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5782] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 5783] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5784] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5785] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 5786] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 5787] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 5788] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5789] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5790] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 5791] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 5792] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5793] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 5794] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 5795] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5796] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5797] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 5798] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5799] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 5800] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 5801] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 5802] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 5803] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5804] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 5805] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 5806] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 5807] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 5808] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5809] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5810] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 5811] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5812] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 5813] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 5814] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5815] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[ 5816] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 5817] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5818] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5819] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 5820] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 5821] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 5822] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5823] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 5824] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 5825] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5826] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 5827] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5828] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5829] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5830] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5831] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 5832] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5833] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5834] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5835] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 5836] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 5837] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 5838] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 5839] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5840] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 5841] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 5842] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 5843] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 5844] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 5845] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 5846] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5847] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 5848] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 5849] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5850] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 5851] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5852] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 5853] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 5854] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 5855] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5856] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 5857] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 5858] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5859] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5860] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5861] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5862] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5863] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 5864] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 5865] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5866] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5867] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 5868] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5869] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5870] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5871] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 5872] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5873] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 5874] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 5875] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5876] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 5877] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5878] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5879] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5880] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 5881] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5882] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 5883] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 5884] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 5885] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5886] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 5887] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5888] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 5889] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 5890] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 5891] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 5892] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5893] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5894] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5895] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 5896] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 5897] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 5898] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5899] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5900] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5901] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5902] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5903] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5904] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5905] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 5906] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 5907] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5908] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 5909] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 5910] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5911] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5912] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 5913] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 5914] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5915] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5916] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 5917] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 5918] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5919] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 5920] = 32'b01000010110111000000000000000000;
	assign	noise_gru_input_weights_array[ 5921] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5922] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 5923] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 5924] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5925] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5926] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 5927] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5928] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 5929] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 5930] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 5931] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5932] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5933] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5934] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5935] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 5936] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 5937] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 5938] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 5939] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 5940] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 5941] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 5942] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5943] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 5944] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 5945] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 5946] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 5947] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5948] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 5949] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 5950] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 5951] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 5952] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5953] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 5954] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 5955] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 5956] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5957] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 5958] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 5959] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 5960] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5961] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5962] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 5963] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 5964] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 5965] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 5966] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 5967] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 5968] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 5969] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 5970] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 5971] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5972] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5973] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 5974] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 5975] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 5976] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 5977] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 5978] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 5979] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 5980] = 32'b11000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 5981] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 5982] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5983] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 5984] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 5985] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 5986] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5987] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 5988] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 5989] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 5990] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 5991] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 5992] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 5993] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 5994] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 5995] = 32'b11000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 5996] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 5997] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 5998] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 5999] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 6000] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6001] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6002] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 6003] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6004] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6005] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 6006] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6007] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 6008] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6009] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 6010] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6011] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6012] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 6013] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6014] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 6015] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 6016] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6017] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6018] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6019] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 6020] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6021] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 6022] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6023] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6024] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 6025] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6026] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6027] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 6028] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6029] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 6030] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 6031] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6032] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 6033] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 6034] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6035] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6036] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 6037] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6038] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 6039] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 6040] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6041] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6042] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 6043] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6044] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 6045] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6046] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6047] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 6048] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 6049] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 6050] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6051] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 6052] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6053] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 6054] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 6055] = 32'b01000010110111000000000000000000;
	assign	noise_gru_input_weights_array[ 6056] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 6057] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 6058] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 6059] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 6060] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 6061] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 6062] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 6063] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 6064] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 6065] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6066] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 6067] = 32'b11000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6068] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6069] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 6070] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 6071] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6072] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 6073] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 6074] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6075] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 6076] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 6077] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 6078] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6079] = 32'b01000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6080] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6081] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 6082] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6083] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6084] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6085] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6086] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6087] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 6088] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6089] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6090] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 6091] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6092] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 6093] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6094] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6095] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 6096] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6097] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 6098] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 6099] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 6100] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 6101] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6102] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6103] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 6104] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6105] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6106] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6107] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6108] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6109] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 6110] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 6111] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 6112] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 6113] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 6114] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6115] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6116] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 6117] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 6118] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 6119] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 6120] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 6121] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6122] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6123] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6124] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6125] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6126] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6127] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 6128] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6129] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6130] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 6131] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6132] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 6133] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 6134] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6135] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 6136] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6137] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6138] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 6139] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6140] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 6141] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 6142] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 6143] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6144] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 6145] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 6146] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6147] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 6148] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6149] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 6150] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6151] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 6152] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6153] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6154] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 6155] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 6156] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6157] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 6158] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 6159] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 6160] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 6161] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 6162] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 6163] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 6164] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 6165] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 6166] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 6167] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 6168] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6169] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6170] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 6171] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6172] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 6173] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6174] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 6175] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6176] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 6177] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 6178] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 6179] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 6180] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 6181] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6182] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 6183] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6184] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6185] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 6186] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6187] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6188] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 6189] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 6190] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 6191] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6192] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6193] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 6194] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 6195] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6196] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6197] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 6198] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 6199] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 6200] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 6201] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 6202] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6203] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 6204] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 6205] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 6206] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6207] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6208] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 6209] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 6210] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 6211] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6212] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 6213] = 32'b01000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 6214] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6215] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 6216] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6217] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6218] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 6219] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 6220] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 6221] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6222] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6223] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 6224] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 6225] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 6226] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6227] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 6228] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 6229] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 6230] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6231] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6232] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 6233] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6234] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 6235] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6236] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 6237] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 6238] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6239] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6240] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6241] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 6242] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 6243] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6244] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6245] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 6246] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 6247] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 6248] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 6249] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 6250] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6251] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 6252] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6253] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 6254] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 6255] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6256] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6257] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6258] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6259] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6260] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 6261] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6262] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 6263] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6264] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 6265] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 6266] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6267] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 6268] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6269] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 6270] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6271] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 6272] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6273] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 6274] = 32'b11000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6275] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 6276] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6277] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6278] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6279] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6280] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6281] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6282] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6283] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 6284] = 32'b11000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 6285] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6286] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 6287] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6288] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6289] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6290] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 6291] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6292] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6293] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 6294] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6295] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6296] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 6297] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6298] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6299] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 6300] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 6301] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 6302] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 6303] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6304] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6305] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6306] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 6307] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 6308] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6309] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6310] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6311] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 6312] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6313] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6314] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6315] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6316] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6317] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6318] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 6319] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6320] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 6321] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 6322] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6323] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 6324] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 6325] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6326] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6327] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6328] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6329] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 6330] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6331] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6332] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6333] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 6334] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6335] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6336] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 6337] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 6338] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 6339] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 6340] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 6341] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 6342] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 6343] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6344] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 6345] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6346] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 6347] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 6348] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6349] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6350] = 32'b01000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 6351] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 6352] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 6353] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 6354] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 6355] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6356] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6357] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 6358] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6359] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6360] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 6361] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 6362] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6363] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 6364] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6365] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 6366] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 6367] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 6368] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6369] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6370] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 6371] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6372] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 6373] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6374] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6375] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 6376] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 6377] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6378] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 6379] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 6380] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6381] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6382] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6383] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6384] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6385] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6386] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6387] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 6388] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 6389] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 6390] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 6391] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 6392] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6393] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6394] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 6395] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6396] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 6397] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6398] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 6399] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6400] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6401] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6402] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6403] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6404] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6405] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 6406] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6407] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6408] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 6409] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6410] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 6411] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6412] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 6413] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 6414] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6415] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 6416] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 6417] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6418] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 6419] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 6420] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6421] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6422] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6423] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 6424] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6425] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 6426] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 6427] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 6428] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 6429] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 6430] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6431] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 6432] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6433] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6434] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 6435] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 6436] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6437] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 6438] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6439] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 6440] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 6441] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6442] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6443] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 6444] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6445] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6446] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 6447] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 6448] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 6449] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6450] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6451] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6452] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 6453] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6454] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6455] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 6456] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6457] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 6458] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6459] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6460] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6461] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6462] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6463] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 6464] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 6465] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6466] = 32'b11000010110010100000000000000000;
	assign	noise_gru_input_weights_array[ 6467] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 6468] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6469] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 6470] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6471] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 6472] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6473] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6474] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 6475] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6476] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 6477] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 6478] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6479] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6480] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 6481] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6482] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 6483] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6484] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6485] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 6486] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 6487] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 6488] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6489] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 6490] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 6491] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 6492] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 6493] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 6494] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6495] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6496] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 6497] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 6498] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6499] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6500] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 6501] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6502] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 6503] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6504] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 6505] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 6506] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6507] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 6508] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 6509] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6510] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 6511] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6512] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 6513] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6514] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 6515] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 6516] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 6517] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 6518] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 6519] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6520] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 6521] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 6522] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6523] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 6524] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6525] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6526] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 6527] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 6528] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 6529] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 6530] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6531] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 6532] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6533] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 6534] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6535] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 6536] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 6537] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6538] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 6539] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 6540] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 6541] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 6542] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 6543] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 6544] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 6545] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6546] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6547] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6548] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6549] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 6550] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 6551] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6552] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 6553] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 6554] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 6555] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 6556] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6557] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 6558] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 6559] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6560] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 6561] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 6562] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 6563] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 6564] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6565] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 6566] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 6567] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6568] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 6569] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 6570] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6571] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 6572] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 6573] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6574] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 6575] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6576] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6577] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 6578] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 6579] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6580] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6581] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6582] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6583] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 6584] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 6585] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6586] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 6587] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6588] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 6589] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 6590] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6591] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 6592] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 6593] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6594] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 6595] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6596] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6597] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6598] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 6599] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6600] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 6601] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 6602] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6603] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6604] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 6605] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6606] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 6607] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 6608] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 6609] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6610] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6611] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6612] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6613] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 6614] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 6615] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6616] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 6617] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 6618] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6619] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6620] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 6621] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 6622] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 6623] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6624] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 6625] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6626] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 6627] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 6628] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 6629] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 6630] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 6631] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6632] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6633] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6634] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 6635] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 6636] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 6637] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6638] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 6639] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6640] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6641] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6642] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6643] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 6644] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6645] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6646] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 6647] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6648] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6649] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 6650] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 6651] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 6652] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6653] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 6654] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6655] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 6656] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 6657] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6658] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[ 6659] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 6660] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 6661] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 6662] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 6663] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 6664] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 6665] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 6666] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6667] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 6668] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6669] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 6670] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 6671] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 6672] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 6673] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 6674] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 6675] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6676] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 6677] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6678] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 6679] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6680] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 6681] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 6682] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 6683] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 6684] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 6685] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 6686] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 6687] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 6688] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6689] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6690] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 6691] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 6692] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 6693] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 6694] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 6695] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 6696] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 6697] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 6698] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 6699] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 6700] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 6701] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6702] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6703] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 6704] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 6705] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6706] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6707] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6708] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6709] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6710] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 6711] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6712] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 6713] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 6714] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 6715] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 6716] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 6717] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6718] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6719] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6720] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6721] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 6722] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6723] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 6724] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 6725] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6726] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 6727] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6728] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 6729] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 6730] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6731] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 6732] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 6733] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6734] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6735] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6736] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 6737] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 6738] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 6739] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 6740] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6741] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6742] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6743] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6744] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6745] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6746] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 6747] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 6748] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6749] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6750] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 6751] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6752] = 32'b01000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 6753] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6754] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6755] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 6756] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 6757] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 6758] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 6759] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6760] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 6761] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 6762] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6763] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 6764] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6765] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6766] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 6767] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 6768] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6769] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6770] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6771] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 6772] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6773] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 6774] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 6775] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6776] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6777] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 6778] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 6779] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6780] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6781] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 6782] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 6783] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 6784] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 6785] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 6786] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6787] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 6788] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 6789] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 6790] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6791] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 6792] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 6793] = 32'b11000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 6794] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 6795] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 6796] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6797] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6798] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6799] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 6800] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 6801] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6802] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 6803] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 6804] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 6805] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6806] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 6807] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 6808] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 6809] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 6810] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 6811] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 6812] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6813] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6814] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6815] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 6816] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 6817] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6818] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6819] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6820] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6821] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6822] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6823] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6824] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 6825] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6826] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 6827] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6828] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6829] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6830] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 6831] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 6832] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 6833] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6834] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6835] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 6836] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 6837] = 32'b01000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 6838] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 6839] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6840] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 6841] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 6842] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6843] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6844] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6845] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6846] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 6847] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 6848] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 6849] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 6850] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 6851] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6852] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6853] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 6854] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 6855] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6856] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 6857] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6858] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 6859] = 32'b01000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 6860] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6861] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6862] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6863] = 32'b01000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 6864] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6865] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6866] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6867] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6868] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6869] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 6870] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6871] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 6872] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6873] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 6874] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 6875] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 6876] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6877] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 6878] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 6879] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 6880] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 6881] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 6882] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 6883] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 6884] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6885] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 6886] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 6887] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6888] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 6889] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6890] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6891] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6892] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6893] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 6894] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 6895] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6896] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 6897] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6898] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6899] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6900] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 6901] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6902] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6903] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 6904] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6905] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6906] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6907] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 6908] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 6909] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6910] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 6911] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6912] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6913] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6914] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6915] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6916] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6917] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6918] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 6919] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6920] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6921] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6922] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6923] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6924] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6925] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 6926] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6927] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 6928] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6929] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6930] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6931] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 6932] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 6933] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6934] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6935] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6936] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 6937] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6938] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6939] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6940] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6941] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6942] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6943] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6944] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6945] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 6946] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 6947] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 6948] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6949] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6950] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6951] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 6952] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6953] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6954] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6955] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 6956] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6957] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 6958] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 6959] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6960] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 6961] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6962] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6963] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 6964] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6965] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6966] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 6967] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 6968] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6969] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 6970] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 6971] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6972] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 6973] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 6974] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 6975] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6976] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6977] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6978] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 6979] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6980] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 6981] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 6982] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 6983] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6984] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 6985] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 6986] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 6987] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 6988] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 6989] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6990] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 6991] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 6992] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 6993] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 6994] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 6995] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 6996] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 6997] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 6998] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 6999] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 7000] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7001] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7002] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 7003] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7004] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7005] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7006] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7007] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 7008] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7009] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7010] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7011] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7012] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7013] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 7014] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7015] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7016] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7017] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7018] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7019] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7020] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7021] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 7022] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7023] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 7024] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 7025] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7026] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7027] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7028] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7029] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7030] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7031] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7032] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 7033] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7034] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7035] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7036] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7037] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7038] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7039] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7040] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 7041] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 7042] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7043] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7044] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7045] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7046] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7047] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7048] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7049] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7050] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7051] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7052] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7053] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7054] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7055] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7056] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 7057] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7058] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7059] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 7060] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7061] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7062] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 7063] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 7064] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7065] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7066] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7067] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7068] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7069] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 7070] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7071] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7072] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7073] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7074] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 7075] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7076] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 7077] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7078] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7079] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7080] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7081] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7082] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7083] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7084] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 7085] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7086] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7087] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 7088] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7089] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7090] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7091] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7092] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7093] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 7094] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 7095] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7096] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 7097] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 7098] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 7099] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7100] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7101] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7102] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 7103] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7104] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 7105] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7106] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 7107] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 7108] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7109] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7110] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 7111] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 7112] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 7113] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 7114] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 7115] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7116] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7117] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 7118] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7119] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 7120] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7121] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 7122] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 7123] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 7124] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7125] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7126] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 7127] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 7128] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 7129] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7130] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 7131] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 7132] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7133] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7134] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 7135] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 7136] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 7137] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 7138] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 7139] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7140] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7141] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7142] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 7143] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 7144] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7145] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7146] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7147] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7148] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 7149] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7150] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7151] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7152] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 7153] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 7154] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 7155] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7156] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7157] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7158] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 7159] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7160] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7161] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 7162] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 7163] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 7164] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7165] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7166] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7167] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 7168] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 7169] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7170] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 7171] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 7172] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7173] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 7174] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7175] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 7176] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7177] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7178] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 7179] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7180] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 7181] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7182] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 7183] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7184] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 7185] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 7186] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7187] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7188] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7189] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7190] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7191] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7192] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 7193] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7194] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7195] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7196] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 7197] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 7198] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 7199] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 7200] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 7201] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 7202] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 7203] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 7204] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7205] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 7206] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7207] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 7208] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7209] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7210] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 7211] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7212] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7213] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7214] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 7215] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7216] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7217] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 7218] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7219] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7220] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 7221] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7222] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 7223] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7224] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7225] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7226] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7227] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 7228] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 7229] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 7230] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7231] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 7232] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7233] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7234] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7235] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7236] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 7237] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 7238] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7239] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 7240] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7241] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 7242] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7243] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7244] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7245] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7246] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 7247] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 7248] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 7249] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7250] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 7251] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7252] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7253] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 7254] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7255] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7256] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 7257] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 7258] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 7259] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7260] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7261] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7262] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 7263] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 7264] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7265] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 7266] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7267] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[ 7268] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7269] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7270] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 7271] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 7272] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 7273] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 7274] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7275] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 7276] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7277] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7278] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 7279] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 7280] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 7281] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7282] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7283] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 7284] = 32'b01000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7285] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 7286] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7287] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 7288] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 7289] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 7290] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 7291] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7292] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7293] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7294] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 7295] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 7296] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7297] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7298] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7299] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7300] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 7301] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 7302] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 7303] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 7304] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 7305] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[ 7306] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 7307] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7308] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7309] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7310] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7311] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7312] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 7313] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7314] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7315] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7316] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7317] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 7318] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7319] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 7320] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 7321] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7322] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7323] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 7324] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7325] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7326] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 7327] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7328] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7329] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 7330] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7331] = 32'b11000010110111000000000000000000;
	assign	noise_gru_input_weights_array[ 7332] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 7333] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7334] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7335] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 7336] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 7337] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7338] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7339] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 7340] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7341] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7342] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 7343] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 7344] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 7345] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 7346] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 7347] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7348] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7349] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7350] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 7351] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 7352] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7353] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7354] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7355] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7356] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7357] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7358] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 7359] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7360] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7361] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 7362] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 7363] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 7364] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 7365] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7366] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 7367] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7368] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7369] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7370] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 7371] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7372] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7373] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7374] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 7375] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 7376] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 7377] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 7378] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7379] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 7380] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 7381] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 7382] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7383] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7384] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7385] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 7386] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 7387] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7388] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7389] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7390] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 7391] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7392] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 7393] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7394] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 7395] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7396] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7397] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 7398] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 7399] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7400] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7401] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 7402] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7403] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7404] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7405] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7406] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 7407] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7408] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7409] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 7410] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 7411] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7412] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7413] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 7414] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7415] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 7416] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 7417] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 7418] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7419] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 7420] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 7421] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7422] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7423] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 7424] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7425] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 7426] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7427] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7428] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 7429] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 7430] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 7431] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7432] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 7433] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 7434] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7435] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 7436] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7437] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7438] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 7439] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 7440] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 7441] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 7442] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7443] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7444] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7445] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 7446] = 32'b11000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 7447] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 7448] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7449] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 7450] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7451] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7452] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 7453] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 7454] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 7455] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7456] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7457] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7458] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7459] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 7460] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 7461] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 7462] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 7463] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7464] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 7465] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7466] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 7467] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 7468] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7469] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7470] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7471] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7472] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7473] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7474] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 7475] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 7476] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7477] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 7478] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 7479] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 7480] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 7481] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7482] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7483] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7484] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7485] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 7486] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7487] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 7488] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 7489] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7490] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 7491] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7492] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7493] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7494] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7495] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7496] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7497] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7498] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7499] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 7500] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7501] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7502] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 7503] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7504] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7505] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7506] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7507] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7508] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 7509] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 7510] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7511] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7512] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 7513] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7514] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 7515] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7516] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 7517] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7518] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 7519] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 7520] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7521] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7522] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7523] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 7524] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7525] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 7526] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7527] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 7528] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 7529] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7530] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 7531] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 7532] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7533] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7534] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 7535] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 7536] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 7537] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 7538] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 7539] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 7540] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 7541] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 7542] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7543] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 7544] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7545] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7546] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 7547] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 7548] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7549] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 7550] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 7551] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 7552] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 7553] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 7554] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7555] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 7556] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7557] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 7558] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7559] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 7560] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 7561] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 7562] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7563] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 7564] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7565] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 7566] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 7567] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 7568] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7569] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7570] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7571] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 7572] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 7573] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7574] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7575] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7576] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7577] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 7578] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7579] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7580] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 7581] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7582] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 7583] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 7584] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 7585] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 7586] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7587] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7588] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7589] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 7590] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7591] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 7592] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 7593] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 7594] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 7595] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7596] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7597] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7598] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7599] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7600] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7601] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7602] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7603] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7604] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7605] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 7606] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7607] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 7608] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7609] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7610] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 7611] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 7612] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 7613] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7614] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 7615] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 7616] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7617] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 7618] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 7619] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 7620] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7621] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7622] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 7623] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7624] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 7625] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7626] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7627] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7628] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7629] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 7630] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 7631] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7632] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 7633] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 7634] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7635] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 7636] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7637] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7638] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 7639] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 7640] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7641] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7642] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7643] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7644] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7645] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7646] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7647] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7648] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 7649] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7650] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7651] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 7652] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7653] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7654] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7655] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7656] = 32'b01000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 7657] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 7658] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7659] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 7660] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 7661] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7662] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7663] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7664] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 7665] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 7666] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 7667] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7668] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7669] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 7670] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7671] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 7672] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7673] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 7674] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 7675] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7676] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 7677] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 7678] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7679] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 7680] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 7681] = 32'b01000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7682] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7683] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7684] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 7685] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7686] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 7687] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 7688] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 7689] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 7690] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 7691] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 7692] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7693] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7694] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 7695] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 7696] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7697] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 7698] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7699] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7700] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7701] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 7702] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 7703] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 7704] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 7705] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 7706] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7707] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 7708] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7709] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7710] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7711] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 7712] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 7713] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7714] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7715] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7716] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7717] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 7718] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 7719] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 7720] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7721] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 7722] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 7723] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7724] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 7725] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 7726] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7727] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 7728] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7729] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 7730] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7731] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7732] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7733] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 7734] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 7735] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7736] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7737] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7738] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 7739] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 7740] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 7741] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7742] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7743] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7744] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 7745] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 7746] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7747] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7748] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7749] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 7750] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7751] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7752] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 7753] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7754] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 7755] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7756] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 7757] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7758] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7759] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7760] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 7761] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 7762] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7763] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 7764] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7765] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7766] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 7767] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 7768] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 7769] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 7770] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 7771] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7772] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 7773] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7774] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7775] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7776] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 7777] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 7778] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 7779] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 7780] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7781] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7782] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 7783] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 7784] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 7785] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 7786] = 32'b11000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 7787] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 7788] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 7789] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 7790] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 7791] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7792] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 7793] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 7794] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7795] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 7796] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 7797] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 7798] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 7799] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7800] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 7801] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 7802] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7803] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7804] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 7805] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 7806] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 7807] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 7808] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 7809] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 7810] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7811] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 7812] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 7813] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 7814] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7815] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 7816] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 7817] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 7818] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 7819] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 7820] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 7821] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7822] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 7823] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 7824] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 7825] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7826] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 7827] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7828] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7829] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7830] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 7831] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 7832] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 7833] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7834] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7835] = 32'b01000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 7836] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 7837] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 7838] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 7839] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 7840] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 7841] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7842] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7843] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7844] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7845] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 7846] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 7847] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 7848] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7849] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 7850] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 7851] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 7852] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 7853] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7854] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 7855] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7856] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7857] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 7858] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 7859] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 7860] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 7861] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 7862] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 7863] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 7864] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 7865] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 7866] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7867] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 7868] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 7869] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 7870] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 7871] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 7872] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7873] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 7874] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 7875] = 32'b01000010110111000000000000000000;
	assign	noise_gru_input_weights_array[ 7876] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 7877] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 7878] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 7879] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7880] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 7881] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 7882] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 7883] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7884] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7885] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7886] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 7887] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 7888] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 7889] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 7890] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 7891] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 7892] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 7893] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 7894] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7895] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 7896] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 7897] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7898] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 7899] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 7900] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 7901] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 7902] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 7903] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 7904] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 7905] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 7906] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 7907] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7908] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 7909] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7910] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 7911] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7912] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 7913] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7914] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 7915] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7916] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 7917] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 7918] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 7919] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7920] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 7921] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7922] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 7923] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 7924] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7925] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7926] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7927] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 7928] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 7929] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7930] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 7931] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7932] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 7933] = 32'b01000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 7934] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 7935] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 7936] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7937] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 7938] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 7939] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7940] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 7941] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 7942] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 7943] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 7944] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7945] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 7946] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 7947] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 7948] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 7949] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7950] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7951] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 7952] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 7953] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 7954] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 7955] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 7956] = 32'b01000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 7957] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 7958] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7959] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 7960] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 7961] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 7962] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 7963] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 7964] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 7965] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 7966] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 7967] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 7968] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7969] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 7970] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 7971] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 7972] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 7973] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 7974] = 32'b01000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 7975] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7976] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 7977] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7978] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 7979] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 7980] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 7981] = 32'b01000010110111000000000000000000;
	assign	noise_gru_input_weights_array[ 7982] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 7983] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 7984] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 7985] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 7986] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 7987] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 7988] = 32'b01000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 7989] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 7990] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 7991] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 7992] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 7993] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 7994] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 7995] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 7996] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 7997] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 7998] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 7999] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 8000] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8001] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 8002] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 8003] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 8004] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8005] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 8006] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 8007] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 8008] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 8009] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 8010] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 8011] = 32'b11000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 8012] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 8013] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8014] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 8015] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 8016] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 8017] = 32'b01000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 8018] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 8019] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 8020] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 8021] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8022] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 8023] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8024] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8025] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8026] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 8027] = 32'b11000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 8028] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 8029] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 8030] = 32'b01000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 8031] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8032] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 8033] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 8034] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 8035] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8036] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8037] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 8038] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8039] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8040] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 8041] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 8042] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8043] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 8044] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 8045] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 8046] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 8047] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8048] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8049] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 8050] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8051] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 8052] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 8053] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 8054] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 8055] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8056] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8057] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8058] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8059] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8060] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 8061] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 8062] = 32'b01000010111001100000000000000000;
	assign	noise_gru_input_weights_array[ 8063] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 8064] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 8065] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 8066] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 8067] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8068] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 8069] = 32'b01000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 8070] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8071] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 8072] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 8073] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 8074] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 8075] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 8076] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 8077] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 8078] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 8079] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8080] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 8081] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8082] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 8083] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 8084] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 8085] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8086] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8087] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 8088] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 8089] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8090] = 32'b01000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 8091] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8092] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 8093] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 8094] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 8095] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 8096] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 8097] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 8098] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8099] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 8100] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 8101] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 8102] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 8103] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8104] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 8105] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8106] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 8107] = 32'b01000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 8108] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 8109] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8110] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8111] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8112] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 8113] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8114] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8115] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8116] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8117] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 8118] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8119] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 8120] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8121] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 8122] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 8123] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 8124] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 8125] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 8126] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 8127] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 8128] = 32'b01000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 8129] = 32'b11000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 8130] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 8131] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8132] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8133] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8134] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 8135] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 8136] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 8137] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 8138] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8139] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 8140] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 8141] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 8142] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 8143] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 8144] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 8145] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 8146] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 8147] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 8148] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8149] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 8150] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 8151] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 8152] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 8153] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 8154] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 8155] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8156] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 8157] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 8158] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 8159] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 8160] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8161] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8162] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 8163] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8164] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 8165] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 8166] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 8167] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8168] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 8169] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8170] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 8171] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8172] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 8173] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8174] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8175] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 8176] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8177] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 8178] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8179] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8180] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 8181] = 32'b11000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 8182] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 8183] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 8184] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 8185] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8186] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8187] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 8188] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8189] = 32'b11000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 8190] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 8191] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 8192] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 8193] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 8194] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 8195] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 8196] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 8197] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 8198] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 8199] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8200] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 8201] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8202] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 8203] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 8204] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 8205] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 8206] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 8207] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8208] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 8209] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 8210] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 8211] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 8212] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8213] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8214] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 8215] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8216] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 8217] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 8218] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 8219] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 8220] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 8221] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 8222] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 8223] = 32'b11000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 8224] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 8225] = 32'b01000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 8226] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 8227] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8228] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 8229] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 8230] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 8231] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 8232] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8233] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 8234] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 8235] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 8236] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8237] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8238] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 8239] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 8240] = 32'b01000010110111000000000000000000;
	assign	noise_gru_input_weights_array[ 8241] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 8242] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 8243] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8244] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 8245] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 8246] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 8247] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 8248] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 8249] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 8250] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 8251] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8252] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 8253] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 8254] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 8255] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 8256] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 8257] = 32'b11000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 8258] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 8259] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 8260] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 8261] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8262] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 8263] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 8264] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 8265] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 8266] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 8267] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 8268] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8269] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8270] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 8271] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 8272] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8273] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8274] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 8275] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 8276] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 8277] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8278] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 8279] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 8280] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 8281] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8282] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 8283] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8284] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 8285] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8286] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8287] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8288] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 8289] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 8290] = 32'b11000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 8291] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 8292] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 8293] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 8294] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 8295] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8296] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8297] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8298] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 8299] = 32'b11000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 8300] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 8301] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 8302] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 8303] = 32'b11000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 8304] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 8305] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 8306] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8307] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 8308] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8309] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8310] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 8311] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8312] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 8313] = 32'b01000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 8314] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 8315] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 8316] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 8317] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 8318] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 8319] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 8320] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 8321] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 8322] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 8323] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 8324] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 8325] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 8326] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 8327] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 8328] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8329] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 8330] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 8331] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 8332] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 8333] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 8334] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8335] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 8336] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 8337] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8338] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 8339] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 8340] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8341] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8342] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8343] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 8344] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 8345] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 8346] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 8347] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 8348] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 8349] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 8350] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 8351] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8352] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 8353] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8354] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8355] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8356] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 8357] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8358] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 8359] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 8360] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8361] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8362] = 32'b01000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 8363] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 8364] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 8365] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 8366] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 8367] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 8368] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 8369] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8370] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 8371] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8372] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 8373] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 8374] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 8375] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 8376] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 8377] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 8378] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 8379] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 8380] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8381] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 8382] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8383] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 8384] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 8385] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 8386] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 8387] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 8388] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 8389] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8390] = 32'b01000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 8391] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8392] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 8393] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 8394] = 32'b11000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 8395] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 8396] = 32'b11000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 8397] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 8398] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 8399] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 8400] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 8401] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8402] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 8403] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 8404] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8405] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 8406] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8407] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8408] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 8409] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8410] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 8411] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 8412] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8413] = 32'b11000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 8414] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 8415] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 8416] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 8417] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 8418] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 8419] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 8420] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 8421] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 8422] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 8423] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 8424] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 8425] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 8426] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 8427] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 8428] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 8429] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 8430] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 8431] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8432] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 8433] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8434] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 8435] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8436] = 32'b01000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 8437] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8438] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 8439] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 8440] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8441] = 32'b11000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 8442] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8443] = 32'b11000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 8444] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 8445] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8446] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 8447] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8448] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 8449] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8450] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8451] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8452] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8453] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 8454] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8455] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8456] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8457] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 8458] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 8459] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 8460] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 8461] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 8462] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 8463] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 8464] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8465] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8466] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8467] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8468] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8469] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8470] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8471] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8472] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8473] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8474] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 8475] = 32'b01000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 8476] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 8477] = 32'b01000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 8478] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 8479] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 8480] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8481] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 8482] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 8483] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 8484] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 8485] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 8486] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 8487] = 32'b11000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 8488] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8489] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 8490] = 32'b11000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 8491] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8492] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 8493] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 8494] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 8495] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8496] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 8497] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 8498] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 8499] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 8500] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 8501] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8502] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 8503] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 8504] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8505] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8506] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8507] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 8508] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 8509] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 8510] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 8511] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 8512] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 8513] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8514] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 8515] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8516] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8517] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 8518] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8519] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 8520] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 8521] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8522] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 8523] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 8524] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8525] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8526] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 8527] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 8528] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 8529] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 8530] = 32'b01000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 8531] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 8532] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8533] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 8534] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 8535] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 8536] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8537] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8538] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 8539] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8540] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 8541] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8542] = 32'b11000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 8543] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 8544] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8545] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 8546] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 8547] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 8548] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 8549] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 8550] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 8551] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 8552] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8553] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 8554] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 8555] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8556] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 8557] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8558] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 8559] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 8560] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 8561] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8562] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 8563] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 8564] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 8565] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8566] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 8567] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8568] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8569] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8570] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 8571] = 32'b01000010111001100000000000000000;
	assign	noise_gru_input_weights_array[ 8572] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 8573] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 8574] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 8575] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 8576] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 8577] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 8578] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 8579] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 8580] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 8581] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 8582] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 8583] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8584] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 8585] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 8586] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 8587] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8588] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 8589] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 8590] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 8591] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8592] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 8593] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8594] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 8595] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 8596] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 8597] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8598] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 8599] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 8600] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8601] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8602] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 8603] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 8604] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8605] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 8606] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8607] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8608] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8609] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 8610] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 8611] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8612] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8613] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8614] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 8615] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8616] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 8617] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 8618] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 8619] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 8620] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 8621] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 8622] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 8623] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 8624] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 8625] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 8626] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 8627] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 8628] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 8629] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 8630] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 8631] = 32'b11000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 8632] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8633] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8634] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 8635] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8636] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 8637] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 8638] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8639] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 8640] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 8641] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 8642] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 8643] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 8644] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 8645] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8646] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8647] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8648] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8649] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8650] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 8651] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 8652] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 8653] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 8654] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 8655] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 8656] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8657] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8658] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 8659] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 8660] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8661] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 8662] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 8663] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 8664] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 8665] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 8666] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8667] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 8668] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 8669] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 8670] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 8671] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 8672] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 8673] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[ 8674] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 8675] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 8676] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 8677] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 8678] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 8679] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 8680] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 8681] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 8682] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 8683] = 32'b01000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 8684] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 8685] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 8686] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 8687] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 8688] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 8689] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 8690] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 8691] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 8692] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8693] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 8694] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 8695] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 8696] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8697] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8698] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 8699] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 8700] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 8701] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 8702] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 8703] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8704] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 8705] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 8706] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 8707] = 32'b01000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 8708] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 8709] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8710] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 8711] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 8712] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 8713] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8714] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 8715] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8716] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8717] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 8718] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 8719] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 8720] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8721] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 8722] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 8723] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 8724] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 8725] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 8726] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 8727] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8728] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8729] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 8730] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 8731] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 8732] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8733] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8734] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8735] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 8736] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 8737] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8738] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 8739] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 8740] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8741] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 8742] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8743] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8744] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 8745] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 8746] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 8747] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8748] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 8749] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 8750] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 8751] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 8752] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 8753] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 8754] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 8755] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8756] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 8757] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8758] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8759] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 8760] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 8761] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 8762] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 8763] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 8764] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8765] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8766] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 8767] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 8768] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 8769] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 8770] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 8771] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 8772] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 8773] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 8774] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 8775] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 8776] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 8777] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 8778] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8779] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 8780] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8781] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 8782] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 8783] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 8784] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8785] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 8786] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 8787] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 8788] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 8789] = 32'b01000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 8790] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 8791] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 8792] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 8793] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 8794] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 8795] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 8796] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 8797] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 8798] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8799] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8800] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 8801] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8802] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 8803] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8804] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 8805] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8806] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8807] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8808] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8809] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 8810] = 32'b11000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 8811] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 8812] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8813] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 8814] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 8815] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 8816] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 8817] = 32'b01000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 8818] = 32'b01000010110111000000000000000000;
	assign	noise_gru_input_weights_array[ 8819] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 8820] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 8821] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 8822] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 8823] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 8824] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 8825] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 8826] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 8827] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 8828] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8829] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 8830] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 8831] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 8832] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 8833] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8834] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8835] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 8836] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8837] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 8838] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 8839] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8840] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8841] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 8842] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 8843] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 8844] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8845] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 8846] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 8847] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 8848] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8849] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 8850] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 8851] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 8852] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 8853] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 8854] = 32'b01000010110111000000000000000000;
	assign	noise_gru_input_weights_array[ 8855] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 8856] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8857] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 8858] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 8859] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 8860] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 8861] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 8862] = 32'b01000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 8863] = 32'b01000010111001100000000000000000;
	assign	noise_gru_input_weights_array[ 8864] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 8865] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 8866] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 8867] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8868] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 8869] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 8870] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8871] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8872] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8873] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 8874] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 8875] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 8876] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 8877] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 8878] = 32'b01000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 8879] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 8880] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8881] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8882] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8883] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 8884] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 8885] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8886] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8887] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8888] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8889] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 8890] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 8891] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8892] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 8893] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 8894] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 8895] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 8896] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 8897] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 8898] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 8899] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8900] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 8901] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 8902] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 8903] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 8904] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 8905] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 8906] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8907] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 8908] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 8909] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8910] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8911] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 8912] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8913] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 8914] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 8915] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 8916] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8917] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8918] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 8919] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8920] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 8921] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 8922] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 8923] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 8924] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 8925] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 8926] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 8927] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 8928] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 8929] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 8930] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 8931] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 8932] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 8933] = 32'b11000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 8934] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 8935] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8936] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8937] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 8938] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8939] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8940] = 32'b11000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 8941] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 8942] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 8943] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 8944] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 8945] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 8946] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 8947] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 8948] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8949] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 8950] = 32'b11000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 8951] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 8952] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 8953] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 8954] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 8955] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8956] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 8957] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 8958] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 8959] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8960] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 8961] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 8962] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 8963] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 8964] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 8965] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 8966] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 8967] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 8968] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 8969] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 8970] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 8971] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 8972] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 8973] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 8974] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 8975] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 8976] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 8977] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 8978] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 8979] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 8980] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 8981] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 8982] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8983] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 8984] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 8985] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 8986] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 8987] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 8988] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 8989] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 8990] = 32'b11000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 8991] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 8992] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 8993] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[ 8994] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 8995] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 8996] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 8997] = 32'b11000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 8998] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 8999] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 9000] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 9001] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 9002] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 9003] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 9004] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9005] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 9006] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 9007] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 9008] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9009] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 9010] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 9011] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 9012] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 9013] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 9014] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 9015] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9016] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 9017] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9018] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9019] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 9020] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 9021] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 9022] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 9023] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 9024] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 9025] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 9026] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 9027] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 9028] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 9029] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 9030] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 9031] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 9032] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 9033] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 9034] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 9035] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 9036] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 9037] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 9038] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9039] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 9040] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 9041] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 9042] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 9043] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 9044] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 9045] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 9046] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 9047] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9048] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 9049] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9050] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9051] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 9052] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9053] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 9054] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9055] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 9056] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 9057] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 9058] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 9059] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 9060] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9061] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 9062] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 9063] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 9064] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 9065] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 9066] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 9067] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 9068] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 9069] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 9070] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 9071] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 9072] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 9073] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 9074] = 32'b11000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 9075] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 9076] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9077] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 9078] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 9079] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9080] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9081] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 9082] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 9083] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 9084] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 9085] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 9086] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 9087] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 9088] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9089] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 9090] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 9091] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 9092] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 9093] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 9094] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9095] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 9096] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 9097] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9098] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 9099] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 9100] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 9101] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 9102] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 9103] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 9104] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 9105] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 9106] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 9107] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 9108] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 9109] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 9110] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 9111] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 9112] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 9113] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 9114] = 32'b11000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 9115] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 9116] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 9117] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9118] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 9119] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9120] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 9121] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 9122] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9123] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 9124] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9125] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 9126] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9127] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 9128] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 9129] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 9130] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 9131] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 9132] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 9133] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[ 9134] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 9135] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 9136] = 32'b01000010111001100000000000000000;
	assign	noise_gru_input_weights_array[ 9137] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 9138] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 9139] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 9140] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 9141] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 9142] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 9143] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 9144] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 9145] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 9146] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 9147] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 9148] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9149] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 9150] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 9151] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 9152] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 9153] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9154] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 9155] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 9156] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 9157] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 9158] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 9159] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 9160] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 9161] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 9162] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9163] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 9164] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 9165] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[ 9166] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 9167] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 9168] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 9169] = 32'b11000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 9170] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9171] = 32'b01000010111001100000000000000000;
	assign	noise_gru_input_weights_array[ 9172] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 9173] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 9174] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 9175] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 9176] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 9177] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 9178] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 9179] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 9180] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 9181] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 9182] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9183] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 9184] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9185] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9186] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 9187] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 9188] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 9189] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9190] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 9191] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 9192] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9193] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 9194] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 9195] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 9196] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9197] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 9198] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 9199] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 9200] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 9201] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9202] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 9203] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9204] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 9205] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 9206] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 9207] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 9208] = 32'b11000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 9209] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 9210] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 9211] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 9212] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 9213] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 9214] = 32'b01000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9215] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9216] = 32'b11000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 9217] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 9218] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9219] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 9220] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 9221] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 9222] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 9223] = 32'b11000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 9224] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 9225] = 32'b01000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 9226] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 9227] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 9228] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 9229] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 9230] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9231] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 9232] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 9233] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9234] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 9235] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9236] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 9237] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9238] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 9239] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9240] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 9241] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 9242] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9243] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 9244] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 9245] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 9246] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9247] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 9248] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 9249] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 9250] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 9251] = 32'b01000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 9252] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 9253] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 9254] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 9255] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 9256] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 9257] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9258] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 9259] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 9260] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 9261] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 9262] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 9263] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 9264] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 9265] = 32'b11000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 9266] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 9267] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9268] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9269] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 9270] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 9271] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 9272] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 9273] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 9274] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 9275] = 32'b11000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 9276] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 9277] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 9278] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 9279] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 9280] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 9281] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9282] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 9283] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 9284] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9285] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 9286] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 9287] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 9288] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9289] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 9290] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 9291] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9292] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9293] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 9294] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 9295] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 9296] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9297] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9298] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 9299] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 9300] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 9301] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 9302] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 9303] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 9304] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9305] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 9306] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 9307] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 9308] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9309] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 9310] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9311] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 9312] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 9313] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9314] = 32'b01000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 9315] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 9316] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 9317] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9318] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 9319] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9320] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 9321] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 9322] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 9323] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9324] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 9325] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9326] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9327] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9328] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 9329] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9330] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 9331] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 9332] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 9333] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 9334] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 9335] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9336] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 9337] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9338] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 9339] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 9340] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9341] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 9342] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9343] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 9344] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 9345] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 9346] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9347] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 9348] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9349] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 9350] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 9351] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9352] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9353] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[ 9354] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9355] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 9356] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 9357] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 9358] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 9359] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9360] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 9361] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 9362] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 9363] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 9364] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 9365] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 9366] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 9367] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 9368] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 9369] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 9370] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 9371] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9372] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9373] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 9374] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 9375] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 9376] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 9377] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9378] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 9379] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9380] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 9381] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9382] = 32'b11000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 9383] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 9384] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 9385] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 9386] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[ 9387] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 9388] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 9389] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 9390] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 9391] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 9392] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 9393] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9394] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 9395] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 9396] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[ 9397] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 9398] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 9399] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9400] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 9401] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 9402] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9403] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9404] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 9405] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 9406] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 9407] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 9408] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 9409] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 9410] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 9411] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 9412] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 9413] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 9414] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 9415] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 9416] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 9417] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 9418] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 9419] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 9420] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 9421] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9422] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 9423] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 9424] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 9425] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 9426] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9427] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 9428] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 9429] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 9430] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9431] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9432] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 9433] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9434] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 9435] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 9436] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 9437] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 9438] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9439] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 9440] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 9441] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9442] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 9443] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9444] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 9445] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 9446] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 9447] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9448] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 9449] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 9450] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 9451] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9452] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 9453] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 9454] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 9455] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 9456] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 9457] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 9458] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 9459] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 9460] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 9461] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 9462] = 32'b11000010110111000000000000000000;
	assign	noise_gru_input_weights_array[ 9463] = 32'b11000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 9464] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 9465] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 9466] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 9467] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 9468] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 9469] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 9470] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 9471] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 9472] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 9473] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9474] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 9475] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9476] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9477] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 9478] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9479] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 9480] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 9481] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 9482] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9483] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 9484] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9485] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 9486] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 9487] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 9488] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 9489] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 9490] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 9491] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[ 9492] = 32'b01000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 9493] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 9494] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9495] = 32'b11000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 9496] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 9497] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 9498] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9499] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 9500] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 9501] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 9502] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 9503] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 9504] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9505] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 9506] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9507] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 9508] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 9509] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9510] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 9511] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 9512] = 32'b01000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 9513] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 9514] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 9515] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9516] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 9517] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 9518] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 9519] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 9520] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 9521] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 9522] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 9523] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 9524] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 9525] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 9526] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 9527] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 9528] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 9529] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 9530] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9531] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9532] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 9533] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 9534] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9535] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 9536] = 32'b11000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 9537] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 9538] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9539] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 9540] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9541] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 9542] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 9543] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 9544] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[ 9545] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 9546] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9547] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 9548] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 9549] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 9550] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 9551] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 9552] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9553] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 9554] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 9555] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 9556] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 9557] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[ 9558] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 9559] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 9560] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 9561] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 9562] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 9563] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9564] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 9565] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 9566] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9567] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 9568] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 9569] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 9570] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9571] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 9572] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 9573] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9574] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 9575] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 9576] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 9577] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 9578] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 9579] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9580] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 9581] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 9582] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 9583] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9584] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 9585] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 9586] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 9587] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[ 9588] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 9589] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 9590] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 9591] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 9592] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 9593] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 9594] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 9595] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9596] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 9597] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 9598] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9599] = 32'b01000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 9600] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 9601] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 9602] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 9603] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 9604] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 9605] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9606] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 9607] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 9608] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 9609] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9610] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 9611] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 9612] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[ 9613] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 9614] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 9615] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 9616] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 9617] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 9618] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9619] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9620] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9621] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 9622] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 9623] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 9624] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9625] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 9626] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 9627] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9628] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 9629] = 32'b01000010111001100000000000000000;
	assign	noise_gru_input_weights_array[ 9630] = 32'b01000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 9631] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 9632] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 9633] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 9634] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 9635] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9636] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 9637] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 9638] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 9639] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 9640] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 9641] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 9642] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 9643] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 9644] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 9645] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 9646] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9647] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 9648] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[ 9649] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 9650] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 9651] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 9652] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9653] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 9654] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 9655] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 9656] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 9657] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 9658] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9659] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 9660] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[ 9661] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 9662] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[ 9663] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 9664] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 9665] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 9666] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 9667] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 9668] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 9669] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 9670] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 9671] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 9672] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 9673] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[ 9674] = 32'b01000010110100000000000000000000;
	assign	noise_gru_input_weights_array[ 9675] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 9676] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9677] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9678] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 9679] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 9680] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[ 9681] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[ 9682] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 9683] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 9684] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 9685] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 9686] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 9687] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 9688] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 9689] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 9690] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 9691] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 9692] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 9693] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 9694] = 32'b11000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 9695] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 9696] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 9697] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 9698] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 9699] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 9700] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 9701] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9702] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[ 9703] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[ 9704] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9705] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 9706] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9707] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 9708] = 32'b11000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 9709] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 9710] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 9711] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 9712] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9713] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 9714] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9715] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 9716] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 9717] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 9718] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 9719] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 9720] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9721] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 9722] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 9723] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 9724] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9725] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 9726] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[ 9727] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[ 9728] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 9729] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[ 9730] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 9731] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 9732] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 9733] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9734] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9735] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 9736] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 9737] = 32'b11000010101110000000000000000000;
	assign	noise_gru_input_weights_array[ 9738] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 9739] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9740] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 9741] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 9742] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 9743] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9744] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 9745] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 9746] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 9747] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 9748] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 9749] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 9750] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9751] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 9752] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 9753] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9754] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 9755] = 32'b11000010110111000000000000000000;
	assign	noise_gru_input_weights_array[ 9756] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 9757] = 32'b11000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 9758] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 9759] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9760] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 9761] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 9762] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 9763] = 32'b11000010110111000000000000000000;
	assign	noise_gru_input_weights_array[ 9764] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 9765] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9766] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[ 9767] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 9768] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 9769] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9770] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 9771] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 9772] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 9773] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 9774] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[ 9775] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9776] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 9777] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9778] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 9779] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[ 9780] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 9781] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[ 9782] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 9783] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 9784] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 9785] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9786] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9787] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[ 9788] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 9789] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 9790] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 9791] = 32'b11000010110110000000000000000000;
	assign	noise_gru_input_weights_array[ 9792] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 9793] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[ 9794] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 9795] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[ 9796] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 9797] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 9798] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9799] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 9800] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9801] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 9802] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 9803] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9804] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[ 9805] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[ 9806] = 32'b01000010110111000000000000000000;
	assign	noise_gru_input_weights_array[ 9807] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 9808] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[ 9809] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9810] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 9811] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[ 9812] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 9813] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 9814] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[ 9815] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9816] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 9817] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9818] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 9819] = 32'b11000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 9820] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 9821] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 9822] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9823] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[ 9824] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 9825] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 9826] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[ 9827] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 9828] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 9829] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 9830] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9831] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 9832] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 9833] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 9834] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[ 9835] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[ 9836] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 9837] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 9838] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9839] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 9840] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 9841] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9842] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9843] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 9844] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[ 9845] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 9846] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9847] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 9848] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 9849] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 9850] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 9851] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[ 9852] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[ 9853] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 9854] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 9855] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9856] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[ 9857] = 32'b11000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 9858] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 9859] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 9860] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[ 9861] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 9862] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9863] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[ 9864] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 9865] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[ 9866] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 9867] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[ 9868] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9869] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[ 9870] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 9871] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[ 9872] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 9873] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[ 9874] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[ 9875] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 9876] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 9877] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 9878] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 9879] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 9880] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9881] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 9882] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[ 9883] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 9884] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9885] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 9886] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 9887] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 9888] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 9889] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9890] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 9891] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 9892] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 9893] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[ 9894] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 9895] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[ 9896] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[ 9897] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 9898] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9899] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 9900] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 9901] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[ 9902] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[ 9903] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[ 9904] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[ 9905] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 9906] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 9907] = 32'b11000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 9908] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[ 9909] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9910] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[ 9911] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[ 9912] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[ 9913] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[ 9914] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[ 9915] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 9916] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9917] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9918] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9919] = 32'b11000010110101000000000000000000;
	assign	noise_gru_input_weights_array[ 9920] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[ 9921] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 9922] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[ 9923] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[ 9924] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 9925] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[ 9926] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[ 9927] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[ 9928] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[ 9929] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9930] = 32'b11000010110011000000000000000000;
	assign	noise_gru_input_weights_array[ 9931] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9932] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[ 9933] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 9934] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9935] = 32'b01000010110100100000000000000000;
	assign	noise_gru_input_weights_array[ 9936] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[ 9937] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 9938] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9939] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9940] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[ 9941] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[ 9942] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9943] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 9944] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[ 9945] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[ 9946] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 9947] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 9948] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9949] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 9950] = 32'b01000010110101100000000000000000;
	assign	noise_gru_input_weights_array[ 9951] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[ 9952] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[ 9953] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 9954] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9955] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9956] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[ 9957] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[ 9958] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 9959] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[ 9960] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[ 9961] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[ 9962] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[ 9963] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[ 9964] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[ 9965] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[ 9966] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 9967] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[ 9968] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 9969] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9970] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[ 9971] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[ 9972] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 9973] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[ 9974] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[ 9975] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 9976] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[ 9977] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[ 9978] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[ 9979] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 9980] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[ 9981] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[ 9982] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[ 9983] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[ 9984] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[ 9985] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[ 9986] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[ 9987] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[ 9988] = 32'b01000010110010000000000000000000;
	assign	noise_gru_input_weights_array[ 9989] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[ 9990] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[ 9991] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[ 9992] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[ 9993] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[ 9994] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[ 9995] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[ 9996] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[ 9997] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[ 9998] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[ 9999] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10000] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[10001] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[10002] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[10003] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[10004] = 32'b01000010111000000000000000000000;
	assign	noise_gru_input_weights_array[10005] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[10006] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[10007] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[10008] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[10009] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[10010] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[10011] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[10012] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[10013] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[10014] = 32'b01000010110010000000000000000000;
	assign	noise_gru_input_weights_array[10015] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10016] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[10017] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[10018] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[10019] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[10020] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[10021] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[10022] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[10023] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[10024] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10025] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[10026] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[10027] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[10028] = 32'b11000010110110000000000000000000;
	assign	noise_gru_input_weights_array[10029] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[10030] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[10031] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[10032] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[10033] = 32'b11000010110010100000000000000000;
	assign	noise_gru_input_weights_array[10034] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[10035] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[10036] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[10037] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[10038] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[10039] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[10040] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[10041] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[10042] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[10043] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[10044] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[10045] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[10046] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[10047] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[10048] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[10049] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[10050] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[10051] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[10052] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[10053] = 32'b01000010110101100000000000000000;
	assign	noise_gru_input_weights_array[10054] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[10055] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[10056] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[10057] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[10058] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[10059] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[10060] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[10061] = 32'b01000010110000000000000000000000;
	assign	noise_gru_input_weights_array[10062] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[10063] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[10064] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[10065] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[10066] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[10067] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10068] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[10069] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[10070] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[10071] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[10072] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[10073] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[10074] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[10075] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[10076] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[10077] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[10078] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10079] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[10080] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[10081] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[10082] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[10083] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[10084] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[10085] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[10086] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[10087] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[10088] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[10089] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[10090] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[10091] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[10092] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[10093] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[10094] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[10095] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[10096] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[10097] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[10098] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[10099] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[10100] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[10101] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[10102] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[10103] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[10104] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[10105] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[10106] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[10107] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[10108] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[10109] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[10110] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[10111] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[10112] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[10113] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[10114] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[10115] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[10116] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[10117] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[10118] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[10119] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[10120] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[10121] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[10122] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[10123] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[10124] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[10125] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[10126] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[10127] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[10128] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[10129] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[10130] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[10131] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[10132] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10133] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[10134] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[10135] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[10136] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[10137] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[10138] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[10139] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[10140] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[10141] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[10142] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[10143] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[10144] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[10145] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[10146] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[10147] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[10148] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[10149] = 32'b11000010110110100000000000000000;
	assign	noise_gru_input_weights_array[10150] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[10151] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[10152] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[10153] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[10154] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[10155] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10156] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[10157] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[10158] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[10159] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[10160] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[10161] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[10162] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[10163] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[10164] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[10165] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[10166] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[10167] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[10168] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[10169] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[10170] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[10171] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[10172] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[10173] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[10174] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[10175] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[10176] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[10177] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[10178] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[10179] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[10180] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[10181] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[10182] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[10183] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[10184] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[10185] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[10186] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[10187] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[10188] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[10189] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[10190] = 32'b01000010111001100000000000000000;
	assign	noise_gru_input_weights_array[10191] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[10192] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[10193] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[10194] = 32'b01000010110100000000000000000000;
	assign	noise_gru_input_weights_array[10195] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[10196] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[10197] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[10198] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[10199] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[10200] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[10201] = 32'b01000010110111000000000000000000;
	assign	noise_gru_input_weights_array[10202] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[10203] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[10204] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[10205] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[10206] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[10207] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[10208] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[10209] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[10210] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[10211] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10212] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[10213] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[10214] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[10215] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[10216] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10217] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[10218] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[10219] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[10220] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[10221] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[10222] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10223] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[10224] = 32'b01000010101111000000000000000000;
	assign	noise_gru_input_weights_array[10225] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[10226] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[10227] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[10228] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[10229] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[10230] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[10231] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[10232] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[10233] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[10234] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[10235] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[10236] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[10237] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[10238] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[10239] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[10240] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[10241] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[10242] = 32'b11000010101110000000000000000000;
	assign	noise_gru_input_weights_array[10243] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[10244] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[10245] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[10246] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[10247] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[10248] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[10249] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[10250] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[10251] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[10252] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[10253] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[10254] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[10255] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[10256] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[10257] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[10258] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[10259] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[10260] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[10261] = 32'b01000010110100000000000000000000;
	assign	noise_gru_input_weights_array[10262] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[10263] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[10264] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[10265] = 32'b11000010110010100000000000000000;
	assign	noise_gru_input_weights_array[10266] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[10267] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[10268] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[10269] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[10270] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[10271] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[10272] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[10273] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[10274] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[10275] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[10276] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[10277] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[10278] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[10279] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[10280] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[10281] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[10282] = 32'b11000010110110100000000000000000;
	assign	noise_gru_input_weights_array[10283] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[10284] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[10285] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[10286] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[10287] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[10288] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[10289] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[10290] = 32'b11000010110111000000000000000000;
	assign	noise_gru_input_weights_array[10291] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[10292] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[10293] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[10294] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[10295] = 32'b11000010110001100000000000000000;
	assign	noise_gru_input_weights_array[10296] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[10297] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[10298] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[10299] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10300] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[10301] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[10302] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[10303] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10304] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[10305] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[10306] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[10307] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[10308] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[10309] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[10310] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[10311] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[10312] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[10313] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[10314] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[10315] = 32'b11000010110110000000000000000000;
	assign	noise_gru_input_weights_array[10316] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[10317] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[10318] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[10319] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[10320] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[10321] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[10322] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[10323] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[10324] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[10325] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[10326] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[10327] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[10328] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[10329] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[10330] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[10331] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[10332] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10333] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[10334] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[10335] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[10336] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[10337] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[10338] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[10339] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[10340] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[10341] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[10342] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10343] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[10344] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[10345] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10346] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[10347] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[10348] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[10349] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[10350] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[10351] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[10352] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[10353] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[10354] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[10355] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[10356] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[10357] = 32'b01000010110111000000000000000000;
	assign	noise_gru_input_weights_array[10358] = 32'b01000010111001100000000000000000;
	assign	noise_gru_input_weights_array[10359] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[10360] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[10361] = 32'b01000010111000000000000000000000;
	assign	noise_gru_input_weights_array[10362] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[10363] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[10364] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[10365] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[10366] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10367] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[10368] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[10369] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[10370] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[10371] = 32'b11000010110111000000000000000000;
	assign	noise_gru_input_weights_array[10372] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[10373] = 32'b11000010110110000000000000000000;
	assign	noise_gru_input_weights_array[10374] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[10375] = 32'b11000010101110000000000000000000;
	assign	noise_gru_input_weights_array[10376] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10377] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[10378] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[10379] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[10380] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[10381] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[10382] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[10383] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[10384] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[10385] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[10386] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[10387] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[10388] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[10389] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[10390] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[10391] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[10392] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[10393] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[10394] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[10395] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[10396] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[10397] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[10398] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10399] = 32'b11000010101110000000000000000000;
	assign	noise_gru_input_weights_array[10400] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[10401] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[10402] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[10403] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[10404] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[10405] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[10406] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[10407] = 32'b01000010101111000000000000000000;
	assign	noise_gru_input_weights_array[10408] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[10409] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[10410] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[10411] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[10412] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[10413] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[10414] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[10415] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[10416] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[10417] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[10418] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[10419] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[10420] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[10421] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[10422] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10423] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[10424] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[10425] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[10426] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[10427] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[10428] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[10429] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[10430] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[10431] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[10432] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[10433] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[10434] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[10435] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[10436] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[10437] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[10438] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[10439] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[10440] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[10441] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[10442] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[10443] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[10444] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[10445] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[10446] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[10447] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[10448] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[10449] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[10450] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[10451] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[10452] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[10453] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[10454] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[10455] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[10456] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[10457] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[10458] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[10459] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[10460] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[10461] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[10462] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10463] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[10464] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[10465] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[10466] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[10467] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10468] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[10469] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[10470] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[10471] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[10472] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[10473] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[10474] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[10475] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[10476] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[10477] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[10478] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[10479] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[10480] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[10481] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[10482] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[10483] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[10484] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[10485] = 32'b11000010110110100000000000000000;
	assign	noise_gru_input_weights_array[10486] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[10487] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[10488] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[10489] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[10490] = 32'b01000010110000000000000000000000;
	assign	noise_gru_input_weights_array[10491] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[10492] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[10493] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[10494] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[10495] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[10496] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[10497] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[10498] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[10499] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[10500] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[10501] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[10502] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[10503] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[10504] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[10505] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[10506] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[10507] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[10508] = 32'b01000010110100000000000000000000;
	assign	noise_gru_input_weights_array[10509] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[10510] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[10511] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[10512] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[10513] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[10514] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[10515] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10516] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[10517] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[10518] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[10519] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[10520] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[10521] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[10522] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[10523] = 32'b11000010110110000000000000000000;
	assign	noise_gru_input_weights_array[10524] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[10525] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[10526] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[10527] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[10528] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[10529] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[10530] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[10531] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[10532] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10533] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[10534] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[10535] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[10536] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[10537] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[10538] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[10539] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[10540] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[10541] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[10542] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[10543] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[10544] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[10545] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[10546] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[10547] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[10548] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[10549] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[10550] = 32'b11000010111001000000000000000000;
	assign	noise_gru_input_weights_array[10551] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[10552] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[10553] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[10554] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[10555] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[10556] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[10557] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[10558] = 32'b11000010110111000000000000000000;
	assign	noise_gru_input_weights_array[10559] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[10560] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[10561] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[10562] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[10563] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[10564] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[10565] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[10566] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[10567] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[10568] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[10569] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[10570] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[10571] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[10572] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[10573] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[10574] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[10575] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[10576] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10577] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[10578] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[10579] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[10580] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[10581] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[10582] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[10583] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[10584] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[10585] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[10586] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[10587] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[10588] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[10589] = 32'b11000010110110000000000000000000;
	assign	noise_gru_input_weights_array[10590] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[10591] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[10592] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[10593] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[10594] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[10595] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[10596] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[10597] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[10598] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[10599] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[10600] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[10601] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[10602] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[10603] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[10604] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[10605] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[10606] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[10607] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[10608] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[10609] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[10610] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[10611] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[10612] = 32'b11000010110111000000000000000000;
	assign	noise_gru_input_weights_array[10613] = 32'b01000010110100100000000000000000;
	assign	noise_gru_input_weights_array[10614] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[10615] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[10616] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[10617] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[10618] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[10619] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[10620] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[10621] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[10622] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[10623] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[10624] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[10625] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[10626] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[10627] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[10628] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[10629] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[10630] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[10631] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[10632] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[10633] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[10634] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[10635] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[10636] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10637] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10638] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[10639] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[10640] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[10641] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[10642] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[10643] = 32'b11000010110111100000000000000000;
	assign	noise_gru_input_weights_array[10644] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[10645] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[10646] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[10647] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[10648] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[10649] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[10650] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[10651] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[10652] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[10653] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[10654] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[10655] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[10656] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[10657] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[10658] = 32'b01000010111000000000000000000000;
	assign	noise_gru_input_weights_array[10659] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[10660] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[10661] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[10662] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[10663] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[10664] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[10665] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[10666] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[10667] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[10668] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[10669] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[10670] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[10671] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[10672] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[10673] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[10674] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[10675] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[10676] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[10677] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[10678] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[10679] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[10680] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[10681] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[10682] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[10683] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[10684] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[10685] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[10686] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[10687] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[10688] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[10689] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[10690] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[10691] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[10692] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[10693] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[10694] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[10695] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[10696] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[10697] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[10698] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[10699] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[10700] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[10701] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[10702] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[10703] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[10704] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[10705] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[10706] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[10707] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[10708] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[10709] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[10710] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[10711] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[10712] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[10713] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[10714] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[10715] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[10716] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[10717] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[10718] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[10719] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[10720] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[10721] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10722] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[10723] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[10724] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[10725] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[10726] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[10727] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[10728] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[10729] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[10730] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[10731] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[10732] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[10733] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[10734] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[10735] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[10736] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[10737] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[10738] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[10739] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[10740] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[10741] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[10742] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[10743] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[10744] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[10745] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[10746] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[10747] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[10748] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[10749] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[10750] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[10751] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[10752] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10753] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[10754] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[10755] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[10756] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[10757] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[10758] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[10759] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[10760] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[10761] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[10762] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[10763] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[10764] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[10765] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[10766] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[10767] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[10768] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[10769] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10770] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[10771] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[10772] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10773] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[10774] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[10775] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[10776] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[10777] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[10778] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[10779] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[10780] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[10781] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[10782] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[10783] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[10784] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[10785] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[10786] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[10787] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[10788] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[10789] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[10790] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[10791] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[10792] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[10793] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[10794] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[10795] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[10796] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[10797] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[10798] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[10799] = 32'b11000010110101000000000000000000;
	assign	noise_gru_input_weights_array[10800] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[10801] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[10802] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[10803] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[10804] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[10805] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[10806] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[10807] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[10808] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[10809] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[10810] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[10811] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[10812] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[10813] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[10814] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[10815] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[10816] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[10817] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[10818] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[10819] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[10820] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[10821] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[10822] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[10823] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[10824] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[10825] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[10826] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[10827] = 32'b11000010111001000000000000000000;
	assign	noise_gru_input_weights_array[10828] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[10829] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[10830] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[10831] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[10832] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[10833] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[10834] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[10835] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[10836] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[10837] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[10838] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[10839] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[10840] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[10841] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[10842] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[10843] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[10844] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[10845] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[10846] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[10847] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[10848] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[10849] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[10850] = 32'b11000010110111000000000000000000;
	assign	noise_gru_input_weights_array[10851] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[10852] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[10853] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[10854] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[10855] = 32'b11000010110011000000000000000000;
	assign	noise_gru_input_weights_array[10856] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[10857] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[10858] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[10859] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[10860] = 32'b01000010110100100000000000000000;
	assign	noise_gru_input_weights_array[10861] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[10862] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[10863] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[10864] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[10865] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[10866] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[10867] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[10868] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[10869] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[10870] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[10871] = 32'b11000010110011000000000000000000;
	assign	noise_gru_input_weights_array[10872] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[10873] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[10874] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[10875] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[10876] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[10877] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[10878] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[10879] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[10880] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[10881] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[10882] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[10883] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[10884] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[10885] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[10886] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[10887] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[10888] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[10889] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[10890] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[10891] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[10892] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[10893] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[10894] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[10895] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[10896] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[10897] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[10898] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[10899] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[10900] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[10901] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[10902] = 32'b01000010111000000000000000000000;
	assign	noise_gru_input_weights_array[10903] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[10904] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[10905] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[10906] = 32'b01000010111001100000000000000000;
	assign	noise_gru_input_weights_array[10907] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[10908] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[10909] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[10910] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[10911] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[10912] = 32'b11000010110001100000000000000000;
	assign	noise_gru_input_weights_array[10913] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[10914] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[10915] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[10916] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[10917] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[10918] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[10919] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[10920] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[10921] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[10922] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[10923] = 32'b01000010111001100000000000000000;
	assign	noise_gru_input_weights_array[10924] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[10925] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[10926] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[10927] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[10928] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[10929] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[10930] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[10931] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[10932] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[10933] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[10934] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[10935] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[10936] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[10937] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[10938] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[10939] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[10940] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[10941] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[10942] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[10943] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[10944] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[10945] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[10946] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[10947] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[10948] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[10949] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[10950] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[10951] = 32'b11000010110110000000000000000000;
	assign	noise_gru_input_weights_array[10952] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[10953] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[10954] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[10955] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[10956] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[10957] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[10958] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[10959] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[10960] = 32'b01000010111000000000000000000000;
	assign	noise_gru_input_weights_array[10961] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[10962] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[10963] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[10964] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[10965] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[10966] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[10967] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[10968] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[10969] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[10970] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[10971] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[10972] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[10973] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[10974] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[10975] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[10976] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[10977] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[10978] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[10979] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[10980] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[10981] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[10982] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[10983] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[10984] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[10985] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[10986] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[10987] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[10988] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[10989] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[10990] = 32'b01000010110100100000000000000000;
	assign	noise_gru_input_weights_array[10991] = 32'b11000010110001100000000000000000;
	assign	noise_gru_input_weights_array[10992] = 32'b01000010110100000000000000000000;
	assign	noise_gru_input_weights_array[10993] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[10994] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[10995] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[10996] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[10997] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[10998] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[10999] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[11000] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[11001] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[11002] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[11003] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[11004] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[11005] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[11006] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[11007] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[11008] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[11009] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[11010] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[11011] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[11012] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[11013] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[11014] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[11015] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[11016] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[11017] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[11018] = 32'b01000010111001100000000000000000;
	assign	noise_gru_input_weights_array[11019] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[11020] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[11021] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[11022] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[11023] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[11024] = 32'b11000010110001100000000000000000;
	assign	noise_gru_input_weights_array[11025] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[11026] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[11027] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[11028] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[11029] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[11030] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[11031] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[11032] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[11033] = 32'b11000010110111100000000000000000;
	assign	noise_gru_input_weights_array[11034] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[11035] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[11036] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[11037] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[11038] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[11039] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[11040] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[11041] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[11042] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11043] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[11044] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[11045] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[11046] = 32'b11000010110111100000000000000000;
	assign	noise_gru_input_weights_array[11047] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11048] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[11049] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[11050] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[11051] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[11052] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[11053] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[11054] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[11055] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[11056] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[11057] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[11058] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[11059] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[11060] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[11061] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[11062] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[11063] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[11064] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[11065] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[11066] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[11067] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[11068] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[11069] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[11070] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[11071] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[11072] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[11073] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[11074] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[11075] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[11076] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[11077] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[11078] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[11079] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[11080] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[11081] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[11082] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[11083] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[11084] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[11085] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[11086] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[11087] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[11088] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[11089] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[11090] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[11091] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[11092] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[11093] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[11094] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[11095] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[11096] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[11097] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[11098] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[11099] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[11100] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[11101] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[11102] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[11103] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[11104] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[11105] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[11106] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[11107] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[11108] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[11109] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[11110] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[11111] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[11112] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[11113] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[11114] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[11115] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[11116] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[11117] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11118] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[11119] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[11120] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[11121] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[11122] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11123] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[11124] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[11125] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[11126] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[11127] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[11128] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[11129] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[11130] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[11131] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[11132] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[11133] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[11134] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[11135] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[11136] = 32'b01000010110010000000000000000000;
	assign	noise_gru_input_weights_array[11137] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[11138] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[11139] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[11140] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[11141] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[11142] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[11143] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[11144] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[11145] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[11146] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[11147] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[11148] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[11149] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[11150] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[11151] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[11152] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[11153] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[11154] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[11155] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[11156] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[11157] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[11158] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[11159] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[11160] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[11161] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[11162] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[11163] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[11164] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[11165] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[11166] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[11167] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[11168] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[11169] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[11170] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[11171] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[11172] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[11173] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[11174] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[11175] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[11176] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[11177] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[11178] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[11179] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[11180] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[11181] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[11182] = 32'b11000010110111000000000000000000;
	assign	noise_gru_input_weights_array[11183] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[11184] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[11185] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[11186] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[11187] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[11188] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[11189] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[11190] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[11191] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[11192] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[11193] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[11194] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[11195] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[11196] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[11197] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[11198] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[11199] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[11200] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[11201] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[11202] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[11203] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[11204] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[11205] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[11206] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[11207] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[11208] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[11209] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[11210] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[11211] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[11212] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[11213] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11214] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[11215] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[11216] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[11217] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[11218] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[11219] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[11220] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[11221] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[11222] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[11223] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[11224] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[11225] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[11226] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[11227] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[11228] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[11229] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[11230] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[11231] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[11232] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[11233] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[11234] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[11235] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[11236] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[11237] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[11238] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[11239] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[11240] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[11241] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[11242] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[11243] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[11244] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[11245] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[11246] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[11247] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[11248] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[11249] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[11250] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[11251] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[11252] = 32'b11000010110111000000000000000000;
	assign	noise_gru_input_weights_array[11253] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[11254] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[11255] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[11256] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[11257] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[11258] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[11259] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[11260] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[11261] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[11262] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[11263] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11264] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[11265] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[11266] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[11267] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[11268] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[11269] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[11270] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[11271] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[11272] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[11273] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[11274] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[11275] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[11276] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[11277] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[11278] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[11279] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[11280] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[11281] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[11282] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[11283] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[11284] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[11285] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[11286] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[11287] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[11288] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[11289] = 32'b01000010110100000000000000000000;
	assign	noise_gru_input_weights_array[11290] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[11291] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[11292] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[11293] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[11294] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[11295] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[11296] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[11297] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[11298] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[11299] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[11300] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[11301] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[11302] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[11303] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[11304] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[11305] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11306] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[11307] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[11308] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[11309] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[11310] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[11311] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[11312] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[11313] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[11314] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[11315] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[11316] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[11317] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[11318] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[11319] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[11320] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[11321] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[11322] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[11323] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[11324] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[11325] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[11326] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[11327] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[11328] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[11329] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[11330] = 32'b11000010110110100000000000000000;
	assign	noise_gru_input_weights_array[11331] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[11332] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[11333] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[11334] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[11335] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[11336] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[11337] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[11338] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[11339] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[11340] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[11341] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[11342] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[11343] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[11344] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[11345] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[11346] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[11347] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[11348] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[11349] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[11350] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[11351] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[11352] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[11353] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[11354] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[11355] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[11356] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[11357] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11358] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[11359] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[11360] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[11361] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[11362] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[11363] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[11364] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[11365] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[11366] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[11367] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[11368] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[11369] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[11370] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[11371] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[11372] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[11373] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[11374] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[11375] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[11376] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[11377] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[11378] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[11379] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[11380] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[11381] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[11382] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[11383] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[11384] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[11385] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[11386] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[11387] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[11388] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[11389] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[11390] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[11391] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[11392] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[11393] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[11394] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[11395] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[11396] = 32'b11000010110011000000000000000000;
	assign	noise_gru_input_weights_array[11397] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[11398] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[11399] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[11400] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[11401] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[11402] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[11403] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[11404] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[11405] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[11406] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[11407] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[11408] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[11409] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[11410] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[11411] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[11412] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[11413] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[11414] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[11415] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[11416] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[11417] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[11418] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[11419] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[11420] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[11421] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[11422] = 32'b11000010110010100000000000000000;
	assign	noise_gru_input_weights_array[11423] = 32'b01000010111001100000000000000000;
	assign	noise_gru_input_weights_array[11424] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[11425] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[11426] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[11427] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[11428] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[11429] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[11430] = 32'b01000010110100000000000000000000;
	assign	noise_gru_input_weights_array[11431] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[11432] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[11433] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[11434] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[11435] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[11436] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[11437] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[11438] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[11439] = 32'b11000010111001000000000000000000;
	assign	noise_gru_input_weights_array[11440] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[11441] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[11442] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[11443] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[11444] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[11445] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[11446] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[11447] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[11448] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[11449] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[11450] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[11451] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[11452] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[11453] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[11454] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[11455] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[11456] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[11457] = 32'b11000010110111100000000000000000;
	assign	noise_gru_input_weights_array[11458] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[11459] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[11460] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[11461] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[11462] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[11463] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[11464] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[11465] = 32'b01000010111000000000000000000000;
	assign	noise_gru_input_weights_array[11466] = 32'b01000010101100100000000000000000;
	assign	noise_gru_input_weights_array[11467] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[11468] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[11469] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[11470] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[11471] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[11472] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[11473] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[11474] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[11475] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[11476] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[11477] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[11478] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[11479] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[11480] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[11481] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[11482] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[11483] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[11484] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[11485] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[11486] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[11487] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[11488] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[11489] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[11490] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[11491] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[11492] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[11493] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[11494] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[11495] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[11496] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[11497] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[11498] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[11499] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11500] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[11501] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[11502] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[11503] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[11504] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[11505] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[11506] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[11507] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[11508] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[11509] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[11510] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[11511] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[11512] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[11513] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[11514] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[11515] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[11516] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[11517] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[11518] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[11519] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[11520] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[11521] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[11522] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[11523] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[11524] = 32'b01000010110101100000000000000000;
	assign	noise_gru_input_weights_array[11525] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[11526] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[11527] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[11528] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[11529] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[11530] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[11531] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[11532] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[11533] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[11534] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[11535] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[11536] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[11537] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[11538] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[11539] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[11540] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[11541] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[11542] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[11543] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[11544] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[11545] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[11546] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[11547] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[11548] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[11549] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[11550] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[11551] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[11552] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[11553] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[11554] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[11555] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[11556] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[11557] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[11558] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[11559] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[11560] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[11561] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[11562] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[11563] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[11564] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[11565] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[11566] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[11567] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[11568] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[11569] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[11570] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[11571] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[11572] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[11573] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[11574] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[11575] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[11576] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[11577] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[11578] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[11579] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[11580] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[11581] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[11582] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[11583] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[11584] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[11585] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[11586] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[11587] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[11588] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[11589] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[11590] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[11591] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[11592] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[11593] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[11594] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[11595] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[11596] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[11597] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[11598] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[11599] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[11600] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[11601] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[11602] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[11603] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[11604] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[11605] = 32'b01000010101111000000000000000000;
	assign	noise_gru_input_weights_array[11606] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[11607] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[11608] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[11609] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[11610] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11611] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[11612] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[11613] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11614] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[11615] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[11616] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[11617] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[11618] = 32'b01000010110001000000000000000000;
	assign	noise_gru_input_weights_array[11619] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[11620] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[11621] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[11622] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[11623] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[11624] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[11625] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[11626] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[11627] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[11628] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[11629] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[11630] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[11631] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[11632] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[11633] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[11634] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[11635] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[11636] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[11637] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[11638] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[11639] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[11640] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[11641] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[11642] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[11643] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[11644] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[11645] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[11646] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[11647] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[11648] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[11649] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[11650] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[11651] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[11652] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[11653] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[11654] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[11655] = 32'b11000010110011000000000000000000;
	assign	noise_gru_input_weights_array[11656] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[11657] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[11658] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[11659] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[11660] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[11661] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[11662] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[11663] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[11664] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[11665] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[11666] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[11667] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[11668] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[11669] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[11670] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[11671] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[11672] = 32'b11000010111001000000000000000000;
	assign	noise_gru_input_weights_array[11673] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[11674] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[11675] = 32'b11000010110001100000000000000000;
	assign	noise_gru_input_weights_array[11676] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[11677] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[11678] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[11679] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[11680] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[11681] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[11682] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[11683] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[11684] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[11685] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[11686] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[11687] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[11688] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[11689] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[11690] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[11691] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[11692] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[11693] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[11694] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[11695] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[11696] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[11697] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[11698] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[11699] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[11700] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[11701] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[11702] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[11703] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[11704] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[11705] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[11706] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[11707] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[11708] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[11709] = 32'b11000010101101000000000000000000;
	assign	noise_gru_input_weights_array[11710] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[11711] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[11712] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[11713] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[11714] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[11715] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[11716] = 32'b11000010110001100000000000000000;
	assign	noise_gru_input_weights_array[11717] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[11718] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[11719] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[11720] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[11721] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[11722] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[11723] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[11724] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[11725] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[11726] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[11727] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[11728] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[11729] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[11730] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[11731] = 32'b01000010110110000000000000000000;
	assign	noise_gru_input_weights_array[11732] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[11733] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[11734] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[11735] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[11736] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11737] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[11738] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[11739] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[11740] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[11741] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[11742] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[11743] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[11744] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[11745] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[11746] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[11747] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[11748] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[11749] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[11750] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[11751] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[11752] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[11753] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[11754] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[11755] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[11756] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[11757] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[11758] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[11759] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[11760] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[11761] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[11762] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[11763] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[11764] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[11765] = 32'b01000010110111000000000000000000;
	assign	noise_gru_input_weights_array[11766] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[11767] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[11768] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[11769] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[11770] = 32'b11000010110100000000000000000000;
	assign	noise_gru_input_weights_array[11771] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[11772] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[11773] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[11774] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[11775] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[11776] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[11777] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[11778] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[11779] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[11780] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[11781] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[11782] = 32'b11000010110101000000000000000000;
	assign	noise_gru_input_weights_array[11783] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[11784] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[11785] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[11786] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[11787] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[11788] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[11789] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[11790] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[11791] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[11792] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[11793] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[11794] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[11795] = 32'b11000010011010000000000000000000;
	assign	noise_gru_input_weights_array[11796] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[11797] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[11798] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11799] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[11800] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[11801] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[11802] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[11803] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[11804] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[11805] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[11806] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[11807] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[11808] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[11809] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[11810] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[11811] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[11812] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[11813] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[11814] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[11815] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[11816] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11817] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[11818] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[11819] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[11820] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[11821] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[11822] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[11823] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[11824] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[11825] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[11826] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[11827] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[11828] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[11829] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[11830] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[11831] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[11832] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[11833] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[11834] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[11835] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[11836] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[11837] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[11838] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[11839] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[11840] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[11841] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[11842] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[11843] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[11844] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[11845] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[11846] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[11847] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[11848] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[11849] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[11850] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[11851] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[11852] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[11853] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[11854] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[11855] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[11856] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[11857] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[11858] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[11859] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[11860] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[11861] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[11862] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[11863] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[11864] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[11865] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[11866] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[11867] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[11868] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[11869] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[11870] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[11871] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[11872] = 32'b01000010101100000000000000000000;
	assign	noise_gru_input_weights_array[11873] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[11874] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[11875] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[11876] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[11877] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[11878] = 32'b11000010110001100000000000000000;
	assign	noise_gru_input_weights_array[11879] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[11880] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[11881] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[11882] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[11883] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[11884] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11885] = 32'b01000010110101000000000000000000;
	assign	noise_gru_input_weights_array[11886] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[11887] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[11888] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[11889] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[11890] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[11891] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[11892] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[11893] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[11894] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[11895] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[11896] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[11897] = 32'b01000010111000000000000000000000;
	assign	noise_gru_input_weights_array[11898] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[11899] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[11900] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11901] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[11902] = 32'b11000010110111000000000000000000;
	assign	noise_gru_input_weights_array[11903] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[11904] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[11905] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[11906] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[11907] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[11908] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[11909] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[11910] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[11911] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[11912] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11913] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[11914] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[11915] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[11916] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[11917] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[11918] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[11919] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[11920] = 32'b11000010110111100000000000000000;
	assign	noise_gru_input_weights_array[11921] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[11922] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[11923] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[11924] = 32'b11000010110110100000000000000000;
	assign	noise_gru_input_weights_array[11925] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[11926] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[11927] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11928] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[11929] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[11930] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11931] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[11932] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[11933] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[11934] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[11935] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11936] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[11937] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[11938] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[11939] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[11940] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[11941] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[11942] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[11943] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[11944] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[11945] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[11946] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[11947] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[11948] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[11949] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[11950] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[11951] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[11952] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[11953] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[11954] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[11955] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[11956] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[11957] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[11958] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[11959] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[11960] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11961] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[11962] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[11963] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[11964] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[11965] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[11966] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[11967] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[11968] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[11969] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[11970] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[11971] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[11972] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[11973] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[11974] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[11975] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[11976] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[11977] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[11978] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[11979] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[11980] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[11981] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[11982] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[11983] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[11984] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[11985] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[11986] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[11987] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[11988] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[11989] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[11990] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[11991] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[11992] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[11993] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[11994] = 32'b01000010110011100000000000000000;
	assign	noise_gru_input_weights_array[11995] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[11996] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[11997] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[11998] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[11999] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[12000] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[12001] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[12002] = 32'b01000010010101000000000000000000;
	assign	noise_gru_input_weights_array[12003] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[12004] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[12005] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[12006] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[12007] = 32'b01000010101111000000000000000000;
	assign	noise_gru_input_weights_array[12008] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[12009] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[12010] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[12011] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[12012] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[12013] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[12014] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[12015] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[12016] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[12017] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[12018] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[12019] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[12020] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[12021] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[12022] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[12023] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12024] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[12025] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[12026] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[12027] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[12028] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[12029] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[12030] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[12031] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[12032] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[12033] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[12034] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[12035] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[12036] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[12037] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[12038] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[12039] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[12040] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[12041] = 32'b01000010110010000000000000000000;
	assign	noise_gru_input_weights_array[12042] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[12043] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[12044] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[12045] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[12046] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[12047] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[12048] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[12049] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[12050] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[12051] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[12052] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[12053] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[12054] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[12055] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[12056] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[12057] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[12058] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[12059] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[12060] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[12061] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[12062] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[12063] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[12064] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[12065] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[12066] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[12067] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[12068] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[12069] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[12070] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[12071] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12072] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[12073] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[12074] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12075] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[12076] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[12077] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[12078] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[12079] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12080] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[12081] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[12082] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[12083] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[12084] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[12085] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[12086] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[12087] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[12088] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[12089] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[12090] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[12091] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[12092] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[12093] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[12094] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[12095] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[12096] = 32'b11000010101111000000000000000000;
	assign	noise_gru_input_weights_array[12097] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[12098] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[12099] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[12100] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[12101] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[12102] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[12103] = 32'b01000010110100100000000000000000;
	assign	noise_gru_input_weights_array[12104] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12105] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[12106] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[12107] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[12108] = 32'b11000010100101100000000000000000;
	assign	noise_gru_input_weights_array[12109] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[12110] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[12111] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[12112] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[12113] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[12114] = 32'b11000010110001000000000000000000;
	assign	noise_gru_input_weights_array[12115] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[12116] = 32'b01000010110111000000000000000000;
	assign	noise_gru_input_weights_array[12117] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[12118] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12119] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12120] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[12121] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[12122] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[12123] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[12124] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[12125] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[12126] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[12127] = 32'b11000010110001100000000000000000;
	assign	noise_gru_input_weights_array[12128] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[12129] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[12130] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[12131] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[12132] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[12133] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[12134] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[12135] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[12136] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[12137] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[12138] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[12139] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[12140] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[12141] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[12142] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[12143] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[12144] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[12145] = 32'b01000010101010100000000000000000;
	assign	noise_gru_input_weights_array[12146] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[12147] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[12148] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[12149] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[12150] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[12151] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[12152] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[12153] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[12154] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[12155] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[12156] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[12157] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[12158] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[12159] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[12160] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[12161] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[12162] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[12163] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[12164] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[12165] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[12166] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[12167] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[12168] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[12169] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[12170] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[12171] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[12172] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[12173] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[12174] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[12175] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[12176] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[12177] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[12178] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[12179] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[12180] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[12181] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12182] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[12183] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[12184] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[12185] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[12186] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[12187] = 32'b11000010111100100000000000000000;
	assign	noise_gru_input_weights_array[12188] = 32'b01000010111101000000000000000000;
	assign	noise_gru_input_weights_array[12189] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[12190] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[12191] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[12192] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[12193] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[12194] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[12195] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[12196] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[12197] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[12198] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[12199] = 32'b01000010110000000000000000000000;
	assign	noise_gru_input_weights_array[12200] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[12201] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[12202] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[12203] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[12204] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[12205] = 32'b01000010100011100000000000000000;
	assign	noise_gru_input_weights_array[12206] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[12207] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[12208] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[12209] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[12210] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[12211] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[12212] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[12213] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[12214] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[12215] = 32'b11000010110011100000000000000000;
	assign	noise_gru_input_weights_array[12216] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[12217] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[12218] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12219] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[12220] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12221] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[12222] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[12223] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[12224] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[12225] = 32'b01000010111001100000000000000000;
	assign	noise_gru_input_weights_array[12226] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[12227] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12228] = 32'b01000010110000000000000000000000;
	assign	noise_gru_input_weights_array[12229] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[12230] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[12231] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[12232] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[12233] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[12234] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[12235] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[12236] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[12237] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[12238] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[12239] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[12240] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[12241] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[12242] = 32'b01000010011000000000000000000000;
	assign	noise_gru_input_weights_array[12243] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[12244] = 32'b01000010110110100000000000000000;
	assign	noise_gru_input_weights_array[12245] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[12246] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[12247] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[12248] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[12249] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[12250] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[12251] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[12252] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[12253] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[12254] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[12255] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[12256] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[12257] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[12258] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[12259] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[12260] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[12261] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[12262] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[12263] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[12264] = 32'b11000001100100000000000000000000;
	assign	noise_gru_input_weights_array[12265] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[12266] = 32'b01000010111000000000000000000000;
	assign	noise_gru_input_weights_array[12267] = 32'b11000010110110000000000000000000;
	assign	noise_gru_input_weights_array[12268] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[12269] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[12270] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[12271] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[12272] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[12273] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[12274] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[12275] = 32'b01000010101000000000000000000000;
	assign	noise_gru_input_weights_array[12276] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[12277] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[12278] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[12279] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[12280] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[12281] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[12282] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[12283] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[12284] = 32'b11000010111110100000000000000000;
	assign	noise_gru_input_weights_array[12285] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[12286] = 32'b01000010110101100000000000000000;
	assign	noise_gru_input_weights_array[12287] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[12288] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[12289] = 32'b01000010111011100000000000000000;
	assign	noise_gru_input_weights_array[12290] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12291] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[12292] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[12293] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[12294] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[12295] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[12296] = 32'b11000010111001000000000000000000;
	assign	noise_gru_input_weights_array[12297] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[12298] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[12299] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[12300] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[12301] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[12302] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[12303] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[12304] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[12305] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[12306] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[12307] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[12308] = 32'b11000010110110100000000000000000;
	assign	noise_gru_input_weights_array[12309] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[12310] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[12311] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[12312] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[12313] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[12314] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[12315] = 32'b11000010101011100000000000000000;
	assign	noise_gru_input_weights_array[12316] = 32'b01000001101100000000000000000000;
	assign	noise_gru_input_weights_array[12317] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[12318] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[12319] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[12320] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[12321] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[12322] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[12323] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[12324] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[12325] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[12326] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[12327] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[12328] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[12329] = 32'b11000010110101100000000000000000;
	assign	noise_gru_input_weights_array[12330] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[12331] = 32'b01000010110011000000000000000000;
	assign	noise_gru_input_weights_array[12332] = 32'b11000010110111100000000000000000;
	assign	noise_gru_input_weights_array[12333] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[12334] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[12335] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[12336] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[12337] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[12338] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[12339] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[12340] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[12341] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[12342] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[12343] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[12344] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[12345] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[12346] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[12347] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[12348] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[12349] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[12350] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[12351] = 32'b01000010100111100000000000000000;
	assign	noise_gru_input_weights_array[12352] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[12353] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[12354] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[12355] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[12356] = 32'b11000010001010000000000000000000;
	assign	noise_gru_input_weights_array[12357] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[12358] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[12359] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[12360] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[12361] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[12362] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[12363] = 32'b01000010111010100000000000000000;
	assign	noise_gru_input_weights_array[12364] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12365] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12366] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[12367] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[12368] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[12369] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[12370] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[12371] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[12372] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[12373] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[12374] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[12375] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[12376] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[12377] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[12378] = 32'b01000010011100000000000000000000;
	assign	noise_gru_input_weights_array[12379] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[12380] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[12381] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[12382] = 32'b11000010111101000000000000000000;
	assign	noise_gru_input_weights_array[12383] = 32'b01000010110101100000000000000000;
	assign	noise_gru_input_weights_array[12384] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[12385] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[12386] = 32'b01000001111000000000000000000000;
	assign	noise_gru_input_weights_array[12387] = 32'b11000010110110100000000000000000;
	assign	noise_gru_input_weights_array[12388] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[12389] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[12390] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[12391] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[12392] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[12393] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[12394] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[12395] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[12396] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[12397] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[12398] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[12399] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[12400] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[12401] = 32'b11000001111110000000000000000000;
	assign	noise_gru_input_weights_array[12402] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[12403] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[12404] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[12405] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[12406] = 32'b11000010110110100000000000000000;
	assign	noise_gru_input_weights_array[12407] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[12408] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[12409] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[12410] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[12411] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[12412] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[12413] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[12414] = 32'b01000010000100000000000000000000;
	assign	noise_gru_input_weights_array[12415] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[12416] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[12417] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[12418] = 32'b01000010101111100000000000000000;
	assign	noise_gru_input_weights_array[12419] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[12420] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[12421] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[12422] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[12423] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[12424] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12425] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[12426] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12427] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[12428] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[12429] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[12430] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[12431] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[12432] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[12433] = 32'b01000010111000100000000000000000;
	assign	noise_gru_input_weights_array[12434] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[12435] = 32'b11000001101110000000000000000000;
	assign	noise_gru_input_weights_array[12436] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[12437] = 32'b11000010010111000000000000000000;
	assign	noise_gru_input_weights_array[12438] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[12439] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[12440] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12441] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[12442] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[12443] = 32'b01000010111100000000000000000000;
	assign	noise_gru_input_weights_array[12444] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[12445] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[12446] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[12447] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[12448] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[12449] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[12450] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[12451] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[12452] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[12453] = 32'b01000010101011100000000000000000;
	assign	noise_gru_input_weights_array[12454] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[12455] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[12456] = 32'b01000010101101100000000000000000;
	assign	noise_gru_input_weights_array[12457] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[12458] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[12459] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[12460] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[12461] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[12462] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[12463] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12464] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[12465] = 32'b01000010111010000000000000000000;
	assign	noise_gru_input_weights_array[12466] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[12467] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[12468] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[12469] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[12470] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[12471] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[12472] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[12473] = 32'b11000001101010000000000000000000;
	assign	noise_gru_input_weights_array[12474] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[12475] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[12476] = 32'b11000010001101000000000000000000;
	assign	noise_gru_input_weights_array[12477] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[12478] = 32'b11000010110000100000000000000000;
	assign	noise_gru_input_weights_array[12479] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[12480] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[12481] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[12482] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[12483] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[12484] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[12485] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[12486] = 32'b01000010110101100000000000000000;
	assign	noise_gru_input_weights_array[12487] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[12488] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[12489] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12490] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[12491] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[12492] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[12493] = 32'b11000010110111000000000000000000;
	assign	noise_gru_input_weights_array[12494] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[12495] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[12496] = 32'b01000010100001100000000000000000;
	assign	noise_gru_input_weights_array[12497] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[12498] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[12499] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[12500] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[12501] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[12502] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[12503] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[12504] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[12505] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[12506] = 32'b11000010100011100000000000000000;
	assign	noise_gru_input_weights_array[12507] = 32'b01000001110010000000000000000000;
	assign	noise_gru_input_weights_array[12508] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[12509] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[12510] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[12511] = 32'b11000011000000000000000000000000;
	assign	noise_gru_input_weights_array[12512] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[12513] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12514] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[12515] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[12516] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[12517] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[12518] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[12519] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[12520] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[12521] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[12522] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[12523] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[12524] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12525] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[12526] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[12527] = 32'b11000010011111000000000000000000;
	assign	noise_gru_input_weights_array[12528] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[12529] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[12530] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[12531] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[12532] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[12533] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[12534] = 32'b01000010101111000000000000000000;
	assign	noise_gru_input_weights_array[12535] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[12536] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[12537] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[12538] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[12539] = 32'b01000010111011000000000000000000;
	assign	noise_gru_input_weights_array[12540] = 32'b11000010110000000000000000000000;
	assign	noise_gru_input_weights_array[12541] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[12542] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[12543] = 32'b11000010010101000000000000000000;
	assign	noise_gru_input_weights_array[12544] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[12545] = 32'b01000001101010000000000000000000;
	assign	noise_gru_input_weights_array[12546] = 32'b01000010111001100000000000000000;
	assign	noise_gru_input_weights_array[12547] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[12548] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[12549] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[12550] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[12551] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[12552] = 32'b01000010100100100000000000000000;
	assign	noise_gru_input_weights_array[12553] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[12554] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[12555] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[12556] = 32'b11000010101100000000000000000000;
	assign	noise_gru_input_weights_array[12557] = 32'b01000010101111000000000000000000;
	assign	noise_gru_input_weights_array[12558] = 32'b01000001111110000000000000000000;
	assign	noise_gru_input_weights_array[12559] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[12560] = 32'b11000010110001100000000000000000;
	assign	noise_gru_input_weights_array[12561] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[12562] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[12563] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[12564] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[12565] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[12566] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[12567] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[12568] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[12569] = 32'b01000010111001100000000000000000;
	assign	noise_gru_input_weights_array[12570] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[12571] = 32'b11000010111110000000000000000000;
	assign	noise_gru_input_weights_array[12572] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[12573] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[12574] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[12575] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[12576] = 32'b01000010011110000000000000000000;
	assign	noise_gru_input_weights_array[12577] = 32'b11000010010100000000000000000000;
	assign	noise_gru_input_weights_array[12578] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[12579] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[12580] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[12581] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[12582] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[12583] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[12584] = 32'b01000010001100000000000000000000;
	assign	noise_gru_input_weights_array[12585] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[12586] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[12587] = 32'b11000010011011000000000000000000;
	assign	noise_gru_input_weights_array[12588] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[12589] = 32'b01000010110111000000000000000000;
	assign	noise_gru_input_weights_array[12590] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[12591] = 32'b01000010110010000000000000000000;
	assign	noise_gru_input_weights_array[12592] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[12593] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12594] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[12595] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[12596] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12597] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[12598] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[12599] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[12600] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[12601] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[12602] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[12603] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12604] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[12605] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[12606] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[12607] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[12608] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[12609] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[12610] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[12611] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[12612] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[12613] = 32'b01000010010100000000000000000000;
	assign	noise_gru_input_weights_array[12614] = 32'b01000010110111000000000000000000;
	assign	noise_gru_input_weights_array[12615] = 32'b11000010000100000000000000000000;
	assign	noise_gru_input_weights_array[12616] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[12617] = 32'b11000010111000000000000000000000;
	assign	noise_gru_input_weights_array[12618] = 32'b01000010110001100000000000000000;
	assign	noise_gru_input_weights_array[12619] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[12620] = 32'b11000010111000100000000000000000;
	assign	noise_gru_input_weights_array[12621] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[12622] = 32'b11000010010010000000000000000000;
	assign	noise_gru_input_weights_array[12623] = 32'b11000010111001000000000000000000;
	assign	noise_gru_input_weights_array[12624] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[12625] = 32'b11000010011110000000000000000000;
	assign	noise_gru_input_weights_array[12626] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[12627] = 32'b01000010000111000000000000000000;
	assign	noise_gru_input_weights_array[12628] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[12629] = 32'b01000010110111000000000000000000;
	assign	noise_gru_input_weights_array[12630] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[12631] = 32'b11000010110010000000000000000000;
	assign	noise_gru_input_weights_array[12632] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[12633] = 32'b01000010111101100000000000000000;
	assign	noise_gru_input_weights_array[12634] = 32'b01000010111100100000000000000000;
	assign	noise_gru_input_weights_array[12635] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[12636] = 32'b01000010101001000000000000000000;
	assign	noise_gru_input_weights_array[12637] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[12638] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[12639] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[12640] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[12641] = 32'b01000010101010000000000000000000;
	assign	noise_gru_input_weights_array[12642] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[12643] = 32'b11000010101001000000000000000000;
	assign	noise_gru_input_weights_array[12644] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[12645] = 32'b11000010110100100000000000000000;
	assign	noise_gru_input_weights_array[12646] = 32'b01000010110111100000000000000000;
	assign	noise_gru_input_weights_array[12647] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[12648] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[12649] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[12650] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[12651] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[12652] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[12653] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[12654] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[12655] = 32'b11000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12656] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[12657] = 32'b01000010100001000000000000000000;
	assign	noise_gru_input_weights_array[12658] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[12659] = 32'b11000010101010000000000000000000;
	assign	noise_gru_input_weights_array[12660] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[12661] = 32'b11000010000101000000000000000000;
	assign	noise_gru_input_weights_array[12662] = 32'b11000010101101100000000000000000;
	assign	noise_gru_input_weights_array[12663] = 32'b01000001110110000000000000000000;
	assign	noise_gru_input_weights_array[12664] = 32'b01000010101001100000000000000000;
	assign	noise_gru_input_weights_array[12665] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[12666] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[12667] = 32'b01000010101110000000000000000000;
	assign	noise_gru_input_weights_array[12668] = 32'b11000010101000000000000000000000;
	assign	noise_gru_input_weights_array[12669] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[12670] = 32'b01000010100100000000000000000000;
	assign	noise_gru_input_weights_array[12671] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[12672] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[12673] = 32'b01000001100000000000000000000000;
	assign	noise_gru_input_weights_array[12674] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[12675] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[12676] = 32'b11000010110101000000000000000000;
	assign	noise_gru_input_weights_array[12677] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[12678] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[12679] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[12680] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[12681] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[12682] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[12683] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[12684] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[12685] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[12686] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[12687] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[12688] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[12689] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[12690] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[12691] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[12692] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[12693] = 32'b11000010100000000000000000000000;
	assign	noise_gru_input_weights_array[12694] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[12695] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[12696] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[12697] = 32'b01000010011011000000000000000000;
	assign	noise_gru_input_weights_array[12698] = 32'b11000000000000000000000000000000;
	assign	noise_gru_input_weights_array[12699] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[12700] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[12701] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[12702] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[12703] = 32'b11000010100101000000000000000000;
	assign	noise_gru_input_weights_array[12704] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[12705] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[12706] = 32'b01000010000110000000000000000000;
	assign	noise_gru_input_weights_array[12707] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[12708] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[12709] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[12710] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[12711] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[12712] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[12713] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[12714] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[12715] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[12716] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[12717] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[12718] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[12719] = 32'b01000010101110100000000000000000;
	assign	noise_gru_input_weights_array[12720] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[12721] = 32'b01000010001010000000000000000000;
	assign	noise_gru_input_weights_array[12722] = 32'b11000010101110100000000000000000;
	assign	noise_gru_input_weights_array[12723] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[12724] = 32'b11000010001110000000000000000000;
	assign	noise_gru_input_weights_array[12725] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[12726] = 32'b01000001111010000000000000000000;
	assign	noise_gru_input_weights_array[12727] = 32'b01000010010010000000000000000000;
	assign	noise_gru_input_weights_array[12728] = 32'b01000010100111000000000000000000;
	assign	noise_gru_input_weights_array[12729] = 32'b01000010100101100000000000000000;
	assign	noise_gru_input_weights_array[12730] = 32'b01000010011111000000000000000000;
	assign	noise_gru_input_weights_array[12731] = 32'b11000010100100100000000000000000;
	assign	noise_gru_input_weights_array[12732] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[12733] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[12734] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[12735] = 32'b01000010011010000000000000000000;
	assign	noise_gru_input_weights_array[12736] = 32'b11000010101000100000000000000000;
	assign	noise_gru_input_weights_array[12737] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[12738] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[12739] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[12740] = 32'b01000010100010100000000000000000;
	assign	noise_gru_input_weights_array[12741] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[12742] = 32'b11000000110000000000000000000000;
	assign	noise_gru_input_weights_array[12743] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[12744] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[12745] = 32'b11000010001001000000000000000000;
	assign	noise_gru_input_weights_array[12746] = 32'b01000010111110000000000000000000;
	assign	noise_gru_input_weights_array[12747] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[12748] = 32'b01000010001011000000000000000000;
	assign	noise_gru_input_weights_array[12749] = 32'b01000010100000100000000000000000;
	assign	noise_gru_input_weights_array[12750] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[12751] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[12752] = 32'b11000010100111100000000000000000;
	assign	noise_gru_input_weights_array[12753] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[12754] = 32'b01000010001110000000000000000000;
	assign	noise_gru_input_weights_array[12755] = 32'b01000001100010000000000000000000;
	assign	noise_gru_input_weights_array[12756] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[12757] = 32'b11000010011001000000000000000000;
	assign	noise_gru_input_weights_array[12758] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[12759] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[12760] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[12761] = 32'b01000010001000000000000000000000;
	assign	noise_gru_input_weights_array[12762] = 32'b11000010100111000000000000000000;
	assign	noise_gru_input_weights_array[12763] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[12764] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[12765] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[12766] = 32'b11000010101011000000000000000000;
	assign	noise_gru_input_weights_array[12767] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[12768] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[12769] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[12770] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[12771] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[12772] = 32'b01000010111111100000000000000000;
	assign	noise_gru_input_weights_array[12773] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[12774] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[12775] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[12776] = 32'b01000010100010000000000000000000;
	assign	noise_gru_input_weights_array[12777] = 32'b11000010000001000000000000000000;
	assign	noise_gru_input_weights_array[12778] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[12779] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[12780] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[12781] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[12782] = 32'b01000010000001000000000000000000;
	assign	noise_gru_input_weights_array[12783] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[12784] = 32'b11000010010000000000000000000000;
	assign	noise_gru_input_weights_array[12785] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[12786] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[12787] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[12788] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[12789] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[12790] = 32'b01000010110000000000000000000000;
	assign	noise_gru_input_weights_array[12791] = 32'b01000001110100000000000000000000;
	assign	noise_gru_input_weights_array[12792] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[12793] = 32'b01000001110000000000000000000000;
	assign	noise_gru_input_weights_array[12794] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[12795] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[12796] = 32'b01000010010110000000000000000000;
	assign	noise_gru_input_weights_array[12797] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[12798] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[12799] = 32'b11000010111111000000000000000000;
	assign	noise_gru_input_weights_array[12800] = 32'b01000010111111000000000000000000;
	assign	noise_gru_input_weights_array[12801] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[12802] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[12803] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[12804] = 32'b01000000100000000000000000000000;
	assign	noise_gru_input_weights_array[12805] = 32'b11000010100000100000000000000000;
	assign	noise_gru_input_weights_array[12806] = 32'b01000010100101000000000000000000;
	assign	noise_gru_input_weights_array[12807] = 32'b11000010100110100000000000000000;
	assign	noise_gru_input_weights_array[12808] = 32'b11000010000011000000000000000000;
	assign	noise_gru_input_weights_array[12809] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[12810] = 32'b11000000111000000000000000000000;
	assign	noise_gru_input_weights_array[12811] = 32'b11000010100010100000000000000000;
	assign	noise_gru_input_weights_array[12812] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[12813] = 32'b01000001010100000000000000000000;
	assign	noise_gru_input_weights_array[12814] = 32'b00000000000000000000000000000000;
	assign	noise_gru_input_weights_array[12815] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[12816] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[12817] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[12818] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[12819] = 32'b11000010011101000000000000000000;
	assign	noise_gru_input_weights_array[12820] = 32'b01000000110000000000000000000000;
	assign	noise_gru_input_weights_array[12821] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[12822] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[12823] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[12824] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[12825] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[12826] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[12827] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[12828] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[12829] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[12830] = 32'b11000010000010000000000000000000;
	assign	noise_gru_input_weights_array[12831] = 32'b01000001010000000000000000000000;
	assign	noise_gru_input_weights_array[12832] = 32'b11000010001000000000000000000000;
	assign	noise_gru_input_weights_array[12833] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[12834] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[12835] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[12836] = 32'b11000010011100000000000000000000;
	assign	noise_gru_input_weights_array[12837] = 32'b11000010100001000000000000000000;
	assign	noise_gru_input_weights_array[12838] = 32'b01000010110000100000000000000000;
	assign	noise_gru_input_weights_array[12839] = 32'b11000001110110000000000000000000;
	assign	noise_gru_input_weights_array[12840] = 32'b01000010000000000000000000000000;
	assign	noise_gru_input_weights_array[12841] = 32'b01000001101000000000000000000000;
	assign	noise_gru_input_weights_array[12842] = 32'b11000010101111100000000000000000;
	assign	noise_gru_input_weights_array[12843] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[12844] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[12845] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[12846] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[12847] = 32'b01000010011101000000000000000000;
	assign	noise_gru_input_weights_array[12848] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[12849] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[12850] = 32'b01000001000100000000000000000000;
	assign	noise_gru_input_weights_array[12851] = 32'b01000001100100000000000000000000;
	assign	noise_gru_input_weights_array[12852] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[12853] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[12854] = 32'b01000010110100100000000000000000;
	assign	noise_gru_input_weights_array[12855] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[12856] = 32'b01000010001111000000000000000000;
	assign	noise_gru_input_weights_array[12857] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[12858] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[12859] = 32'b01000001001000000000000000000000;
	assign	noise_gru_input_weights_array[12860] = 32'b11000010001111000000000000000000;
	assign	noise_gru_input_weights_array[12861] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[12862] = 32'b01000010111110100000000000000000;
	assign	noise_gru_input_weights_array[12863] = 32'b01000010100110100000000000000000;
	assign	noise_gru_input_weights_array[12864] = 32'b01000010101101000000000000000000;
	assign	noise_gru_input_weights_array[12865] = 32'b01000010000010000000000000000000;
	assign	noise_gru_input_weights_array[12866] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[12867] = 32'b01000010010001000000000000000000;
	assign	noise_gru_input_weights_array[12868] = 32'b01000010100000000000000000000000;
	assign	noise_gru_input_weights_array[12869] = 32'b11000001111000000000000000000000;
	assign	noise_gru_input_weights_array[12870] = 32'b11000010100001100000000000000000;
	assign	noise_gru_input_weights_array[12871] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[12872] = 32'b11000010000000000000000000000000;
	assign	noise_gru_input_weights_array[12873] = 32'b11000001110000000000000000000000;
	assign	noise_gru_input_weights_array[12874] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[12875] = 32'b11000001110010000000000000000000;
	assign	noise_gru_input_weights_array[12876] = 32'b11000010111100000000000000000000;
	assign	noise_gru_input_weights_array[12877] = 32'b00111111100000000000000000000000;
	assign	noise_gru_input_weights_array[12878] = 32'b11000010100010000000000000000000;
	assign	noise_gru_input_weights_array[12879] = 32'b01000010010111000000000000000000;
	assign	noise_gru_input_weights_array[12880] = 32'b01000010101000100000000000000000;
	assign	noise_gru_input_weights_array[12881] = 32'b11000010101010100000000000000000;
	assign	noise_gru_input_weights_array[12882] = 32'b11000001001100000000000000000000;
	assign	noise_gru_input_weights_array[12883] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[12884] = 32'b11000001111010000000000000000000;
	assign	noise_gru_input_weights_array[12885] = 32'b11000010110111000000000000000000;
	assign	noise_gru_input_weights_array[12886] = 32'b01000000000000000000000000000000;
	assign	noise_gru_input_weights_array[12887] = 32'b11000010001100000000000000000000;
	assign	noise_gru_input_weights_array[12888] = 32'b01000010001001000000000000000000;
	assign	noise_gru_input_weights_array[12889] = 32'b11000001010000000000000000000000;
	assign	noise_gru_input_weights_array[12890] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[12891] = 32'b01000000111000000000000000000000;
	assign	noise_gru_input_weights_array[12892] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[12893] = 32'b11000010111011000000000000000000;
	assign	noise_gru_input_weights_array[12894] = 32'b01000010100110000000000000000000;
	assign	noise_gru_input_weights_array[12895] = 32'b11000010100110000000000000000000;
	assign	noise_gru_input_weights_array[12896] = 32'b11000001100010000000000000000000;
	assign	noise_gru_input_weights_array[12897] = 32'b11000010001011000000000000000000;
	assign	noise_gru_input_weights_array[12898] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[12899] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[12900] = 32'b01000010101011000000000000000000;
	assign	noise_gru_input_weights_array[12901] = 32'b11000010111101100000000000000000;
	assign	noise_gru_input_weights_array[12902] = 32'b01000010100011000000000000000000;
	assign	noise_gru_input_weights_array[12903] = 32'b01000010001101000000000000000000;
	assign	noise_gru_input_weights_array[12904] = 32'b11000001010100000000000000000000;
	assign	noise_gru_input_weights_array[12905] = 32'b11000010000111000000000000000000;
	assign	noise_gru_input_weights_array[12906] = 32'b01000010111001000000000000000000;
	assign	noise_gru_input_weights_array[12907] = 32'b11000010100100000000000000000000;
	assign	noise_gru_input_weights_array[12908] = 32'b01000010110010100000000000000000;
	assign	noise_gru_input_weights_array[12909] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[12910] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[12911] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[12912] = 32'b11000010010110000000000000000000;
	assign	noise_gru_input_weights_array[12913] = 32'b11000010010001000000000000000000;
	assign	noise_gru_input_weights_array[12914] = 32'b11000010101110000000000000000000;
	assign	noise_gru_input_weights_array[12915] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[12916] = 32'b11000010111010100000000000000000;
	assign	noise_gru_input_weights_array[12917] = 32'b01000001100110000000000000000000;
	assign	noise_gru_input_weights_array[12918] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[12919] = 32'b11000010111010000000000000000000;
	assign	noise_gru_input_weights_array[12920] = 32'b01000010000101000000000000000000;
	assign	noise_gru_input_weights_array[12921] = 32'b01000001000000000000000000000000;
	assign	noise_gru_input_weights_array[12922] = 32'b01000001011100000000000000000000;
	assign	noise_gru_input_weights_array[12923] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[12924] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[12925] = 32'b11000001101100000000000000000000;
	assign	noise_gru_input_weights_array[12926] = 32'b11000001100000000000000000000000;
	assign	noise_gru_input_weights_array[12927] = 32'b01000001101110000000000000000000;
	assign	noise_gru_input_weights_array[12928] = 32'b11000010101001100000000000000000;
	assign	noise_gru_input_weights_array[12929] = 32'b01000000101000000000000000000000;
	assign	noise_gru_input_weights_array[12930] = 32'b01000010011001000000000000000000;
	assign	noise_gru_input_weights_array[12931] = 32'b01000001011000000000000000000000;
	assign	noise_gru_input_weights_array[12932] = 32'b11000001100110000000000000000000;
	assign	noise_gru_input_weights_array[12933] = 32'b11000001000100000000000000000000;
	assign	noise_gru_input_weights_array[12934] = 32'b01000010010011000000000000000000;
	assign	noise_gru_input_weights_array[12935] = 32'b10111111100000000000000000000000;
	assign	noise_gru_input_weights_array[12936] = 32'b11000001101000000000000000000000;
	assign	noise_gru_input_weights_array[12937] = 32'b11000001110100000000000000000000;
	assign	noise_gru_input_weights_array[12938] = 32'b11000000010000000000000000000000;
	assign	noise_gru_input_weights_array[12939] = 32'b11000001000000000000000000000000;
	assign	noise_gru_input_weights_array[12940] = 32'b01000000010000000000000000000000;
	assign	noise_gru_input_weights_array[12941] = 32'b11000001011000000000000000000000;
	assign	noise_gru_input_weights_array[12942] = 32'b11000010010011000000000000000000;
	assign	noise_gru_input_weights_array[12943] = 32'b01000001001100000000000000000000;
	assign	noise_gru_input_weights_array[12944] = 32'b11000010011000000000000000000000;
	assign	noise_gru_input_weights_array[12945] = 32'b01000001111100000000000000000000;
	assign	noise_gru_input_weights_array[12946] = 32'b11000000101000000000000000000000;
	assign	noise_gru_input_weights_array[12947] = 32'b11000010110110000000000000000000;
	assign	noise_gru_input_weights_array[12948] = 32'b11000001001000000000000000000000;
	assign	noise_gru_input_weights_array[12949] = 32'b11000010111001100000000000000000;
	assign	noise_gru_input_weights_array[12950] = 32'b11000010101100100000000000000000;
	assign	noise_gru_input_weights_array[12951] = 32'b11000010000110000000000000000000;
	assign	noise_gru_input_weights_array[12952] = 32'b11000010100011000000000000000000;
	assign	noise_gru_input_weights_array[12953] = 32'b11000000100000000000000000000000;
	assign	noise_gru_input_weights_array[12954] = 32'b11000001011100000000000000000000;
	assign	noise_gru_input_weights_array[12955] = 32'b11000001111100000000000000000000;
	assign	noise_gru_input_weights_array[12956] = 32'b01000010000011000000000000000000;
	assign	noise_gru_input_weights_array[12957] = 32'b01000010010000000000000000000000;
	assign	noise_gru_input_weights_array[12958] = 32'b11000010111011100000000000000000;
	assign	noise_gru_input_weights_array[12959] = 32'b11000010011111000000000000000000;


	assign	noise_gru_recurrent_weights_array[    0] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[    1] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[    2] = 32'b01000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[    3] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[    4] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[    5] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[    6] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[    7] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[    8] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[    9] = 32'b01000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[   10] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   11] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[   12] = 32'b11000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[   13] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   14] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[   15] = 32'b01000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[   16] = 32'b01000010111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   17] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[   18] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[   19] = 32'b11000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[   20] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[   21] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[   22] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[   23] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[   24] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[   25] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   26] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[   27] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   28] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[   29] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   30] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[   31] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   32] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[   33] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[   34] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   35] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   36] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   37] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[   38] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[   39] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[   40] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[   41] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[   42] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[   43] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   44] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[   45] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[   46] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   47] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[   48] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[   49] = 32'b11000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[   50] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[   51] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[   52] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[   53] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[   54] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[   55] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[   56] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   57] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[   58] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   59] = 32'b01000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[   60] = 32'b01000010110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   61] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[   62] = 32'b01000010110001100000000000000000;
	assign	noise_gru_recurrent_weights_array[   63] = 32'b01000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[   64] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[   65] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   66] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[   67] = 32'b11000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[   68] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[   69] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[   70] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[   71] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[   72] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[   73] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[   74] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   75] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   76] = 32'b11000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[   77] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[   78] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[   79] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[   80] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   81] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[   82] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[   83] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   84] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[   85] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   86] = 32'b11000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[   87] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[   88] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[   89] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[   90] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[   91] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[   92] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   93] = 32'b01000010110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[   94] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[   95] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   96] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[   97] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[   98] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[   99] = 32'b01000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[  100] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  101] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  102] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[  103] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  104] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  105] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  106] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  107] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  108] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  109] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  110] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  111] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  112] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  113] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  114] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  115] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[  116] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  117] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  118] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  119] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  120] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  121] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  122] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  123] = 32'b11000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  124] = 32'b11000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[  125] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  126] = 32'b01000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[  127] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  128] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  129] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  130] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  131] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  132] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  133] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  134] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  135] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  136] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  137] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  138] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  139] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  140] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  141] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  142] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  143] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  144] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  145] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  146] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[  147] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  148] = 32'b01000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[  149] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  150] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  151] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  152] = 32'b11000010111001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  153] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  154] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  155] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  156] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  157] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  158] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  159] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  160] = 32'b01000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  161] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  162] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  163] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[  164] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  165] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  166] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  167] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  168] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  169] = 32'b01000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[  170] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  171] = 32'b01000010110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  172] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  173] = 32'b01000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[  174] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  175] = 32'b01000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  176] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  177] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  178] = 32'b01000010110101100000000000000000;
	assign	noise_gru_recurrent_weights_array[  179] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  180] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  181] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  182] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  183] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  184] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  185] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  186] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  187] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  188] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  189] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  190] = 32'b11000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  191] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  192] = 32'b01000010110001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  193] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  194] = 32'b01000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  195] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  196] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  197] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  198] = 32'b01000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  199] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  200] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  201] = 32'b01000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[  202] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  203] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  204] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  205] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  206] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  207] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  208] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  209] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  210] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  211] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  212] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  213] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  214] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  215] = 32'b11000010110111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  216] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  217] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  218] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  219] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  220] = 32'b11000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[  221] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  222] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  223] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  224] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  225] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  226] = 32'b11000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[  227] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  228] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  229] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  230] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  231] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  232] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  233] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  234] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  235] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  236] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  237] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  238] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  239] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  240] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  241] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  242] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  243] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  244] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  245] = 32'b11000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[  246] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  247] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  248] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  249] = 32'b01000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[  250] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  251] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[  252] = 32'b01000010101100100000000000000000;
	assign	noise_gru_recurrent_weights_array[  253] = 32'b11000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[  254] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  255] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  256] = 32'b11000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[  257] = 32'b11000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[  258] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  259] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  260] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  261] = 32'b11000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[  262] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  263] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  264] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  265] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  266] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  267] = 32'b11000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[  268] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  269] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  270] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  271] = 32'b11000010101110100000000000000000;
	assign	noise_gru_recurrent_weights_array[  272] = 32'b11000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[  273] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  274] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  275] = 32'b01000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[  276] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  277] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  278] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  279] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  280] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  281] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  282] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  283] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  284] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  285] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  286] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  287] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  288] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  289] = 32'b01000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[  290] = 32'b01000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  291] = 32'b01000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[  292] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  293] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  294] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  295] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  296] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  297] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  298] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  299] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  300] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  301] = 32'b01000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[  302] = 32'b01000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[  303] = 32'b01000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[  304] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  305] = 32'b11000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  306] = 32'b01000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  307] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[  308] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  309] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  310] = 32'b11000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[  311] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  312] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  313] = 32'b11000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[  314] = 32'b11000010110101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  315] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  316] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  317] = 32'b01000010110101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  318] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  319] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  320] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  321] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  322] = 32'b01000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[  323] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  324] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[  325] = 32'b01000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[  326] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  327] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  328] = 32'b01000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  329] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[  330] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  331] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  332] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  333] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  334] = 32'b11000010101110100000000000000000;
	assign	noise_gru_recurrent_weights_array[  335] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  336] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  337] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  338] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  339] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  340] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  341] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  342] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  343] = 32'b01000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  344] = 32'b11000010110001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  345] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  346] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[  347] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  348] = 32'b01000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[  349] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  350] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[  351] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  352] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  353] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  354] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  355] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  356] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  357] = 32'b01000010110001100000000000000000;
	assign	noise_gru_recurrent_weights_array[  358] = 32'b11000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[  359] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  360] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  361] = 32'b01000010110001100000000000000000;
	assign	noise_gru_recurrent_weights_array[  362] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  363] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  364] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  365] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  366] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  367] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  368] = 32'b11000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  369] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  370] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  371] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  372] = 32'b01000010111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  373] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  374] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  375] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  376] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  377] = 32'b11000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  378] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  379] = 32'b01000010110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  380] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  381] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  382] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  383] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  384] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  385] = 32'b11000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[  386] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[  387] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  388] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  389] = 32'b11000010111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  390] = 32'b11000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  391] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  392] = 32'b01000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  393] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  394] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  395] = 32'b11000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  396] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  397] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  398] = 32'b11000010111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  399] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  400] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  401] = 32'b01000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[  402] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  403] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[  404] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[  405] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  406] = 32'b01000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  407] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  408] = 32'b11000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  409] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  410] = 32'b01000010110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  411] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  412] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  413] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  414] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  415] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  416] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  417] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  418] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  419] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  420] = 32'b01000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[  421] = 32'b01000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[  422] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  423] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  424] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  425] = 32'b01000010110101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  426] = 32'b11000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  427] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  428] = 32'b01000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  429] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  430] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  431] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  432] = 32'b11000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[  433] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  434] = 32'b01000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[  435] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  436] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  437] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  438] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  439] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  440] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  441] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  442] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  443] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  444] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  445] = 32'b01000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  446] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  447] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  448] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  449] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  450] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  451] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  452] = 32'b01000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[  453] = 32'b11000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[  454] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  455] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  456] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  457] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  458] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  459] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  460] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  461] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  462] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  463] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  464] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  465] = 32'b11000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  466] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  467] = 32'b11000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[  468] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  469] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  470] = 32'b01000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  471] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  472] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  473] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  474] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  475] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  476] = 32'b11000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[  477] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  478] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  479] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  480] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  481] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  482] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  483] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  484] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  485] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  486] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  487] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  488] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  489] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  490] = 32'b11000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[  491] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  492] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  493] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  494] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  495] = 32'b01000010110001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  496] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  497] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  498] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  499] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  500] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  501] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  502] = 32'b11000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  503] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  504] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  505] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  506] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  507] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  508] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  509] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  510] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  511] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  512] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  513] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  514] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  515] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  516] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[  517] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  518] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  519] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  520] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  521] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  522] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[  523] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  524] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  525] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  526] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  527] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  528] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  529] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  530] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[  531] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  532] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  533] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  534] = 32'b11000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  535] = 32'b01000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  536] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  537] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  538] = 32'b11000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  539] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  540] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[  541] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  542] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  543] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  544] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  545] = 32'b11000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[  546] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  547] = 32'b11000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  548] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  549] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  550] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  551] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  552] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  553] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  554] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  555] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  556] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  557] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  558] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  559] = 32'b01000010110111100000000000000000;
	assign	noise_gru_recurrent_weights_array[  560] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  561] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  562] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  563] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  564] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  565] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  566] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  567] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  568] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  569] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  570] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[  571] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  572] = 32'b01000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  573] = 32'b11000010110011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  574] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  575] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  576] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  577] = 32'b01000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[  578] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  579] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  580] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[  581] = 32'b01000010110101100000000000000000;
	assign	noise_gru_recurrent_weights_array[  582] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  583] = 32'b11000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  584] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  585] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  586] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  587] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  588] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  589] = 32'b01000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[  590] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  591] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  592] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  593] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  594] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  595] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  596] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  597] = 32'b11000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  598] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  599] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  600] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  601] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  602] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  603] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  604] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  605] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  606] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  607] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  608] = 32'b11000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  609] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  610] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  611] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  612] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  613] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  614] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  615] = 32'b11000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  616] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  617] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  618] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  619] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  620] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  621] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  622] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  623] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[  624] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  625] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  626] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  627] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  628] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  629] = 32'b01000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  630] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  631] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  632] = 32'b11000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[  633] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  634] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  635] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  636] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  637] = 32'b11000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  638] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  639] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  640] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  641] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[  642] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  643] = 32'b11000010110011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  644] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  645] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  646] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[  647] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  648] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  649] = 32'b11000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  650] = 32'b01000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  651] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  652] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  653] = 32'b01000010110001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  654] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  655] = 32'b01000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[  656] = 32'b11000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[  657] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  658] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  659] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  660] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  661] = 32'b11000010110001100000000000000000;
	assign	noise_gru_recurrent_weights_array[  662] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  663] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  664] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  665] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  666] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  667] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  668] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  669] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  670] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  671] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  672] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  673] = 32'b11000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  674] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  675] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[  676] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  677] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[  678] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  679] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  680] = 32'b01000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  681] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  682] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  683] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  684] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  685] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  686] = 32'b01000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  687] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  688] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  689] = 32'b01000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  690] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  691] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  692] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[  693] = 32'b11000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[  694] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  695] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  696] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  697] = 32'b01000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  698] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  699] = 32'b01000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  700] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  701] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  702] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  703] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  704] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  705] = 32'b01000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[  706] = 32'b11000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[  707] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  708] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  709] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  710] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  711] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  712] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  713] = 32'b01000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  714] = 32'b11000010110001100000000000000000;
	assign	noise_gru_recurrent_weights_array[  715] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  716] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  717] = 32'b01000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  718] = 32'b01000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  719] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  720] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  721] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  722] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  723] = 32'b01000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[  724] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  725] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  726] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  727] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  728] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  729] = 32'b01000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  730] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  731] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  732] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  733] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  734] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  735] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  736] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  737] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  738] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  739] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  740] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  741] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  742] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  743] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  744] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  745] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  746] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  747] = 32'b01000010110101100000000000000000;
	assign	noise_gru_recurrent_weights_array[  748] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  749] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  750] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  751] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  752] = 32'b11000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  753] = 32'b01000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  754] = 32'b01000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  755] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  756] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  757] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  758] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  759] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  760] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  761] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  762] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  763] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  764] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  765] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  766] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  767] = 32'b01000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[  768] = 32'b11000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[  769] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  770] = 32'b01000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[  771] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  772] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  773] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  774] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  775] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  776] = 32'b11000010111001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  777] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  778] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  779] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[  780] = 32'b01000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  781] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  782] = 32'b01000010111001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  783] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  784] = 32'b01000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[  785] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  786] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  787] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  788] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  789] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[  790] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  791] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  792] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  793] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  794] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  795] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  796] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  797] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  798] = 32'b01000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  799] = 32'b11000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  800] = 32'b01000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[  801] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  802] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  803] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  804] = 32'b01000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  805] = 32'b01000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  806] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  807] = 32'b01000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[  808] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  809] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  810] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  811] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  812] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  813] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  814] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  815] = 32'b11000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[  816] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  817] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  818] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  819] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[  820] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  821] = 32'b11000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[  822] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  823] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  824] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  825] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  826] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  827] = 32'b11000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  828] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  829] = 32'b11000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[  830] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  831] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  832] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  833] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  834] = 32'b11000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[  835] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[  836] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  837] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  838] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  839] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  840] = 32'b01000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[  841] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  842] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  843] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  844] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  845] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  846] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  847] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  848] = 32'b01000010110101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  849] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  850] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  851] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  852] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  853] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  854] = 32'b11000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  855] = 32'b11000011000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  856] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  857] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  858] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[  859] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  860] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  861] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  862] = 32'b11000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  863] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[  864] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  865] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  866] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  867] = 32'b11000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  868] = 32'b01000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  869] = 32'b01000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  870] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  871] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  872] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  873] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  874] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  875] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  876] = 32'b01000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[  877] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  878] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  879] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  880] = 32'b11000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  881] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  882] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  883] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[  884] = 32'b11000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  885] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  886] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  887] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  888] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  889] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  890] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  891] = 32'b01000010110001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  892] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  893] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  894] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[  895] = 32'b11000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  896] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  897] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  898] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  899] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  900] = 32'b01000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[  901] = 32'b01000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  902] = 32'b01000010110111100000000000000000;
	assign	noise_gru_recurrent_weights_array[  903] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  904] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  905] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  906] = 32'b11000010110101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  907] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  908] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  909] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  910] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  911] = 32'b01000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[  912] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  913] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  914] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  915] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  916] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  917] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  918] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  919] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  920] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  921] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  922] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  923] = 32'b01000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[  924] = 32'b11000010110111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  925] = 32'b01000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  926] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  927] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  928] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  929] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  930] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  931] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  932] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  933] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  934] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  935] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  936] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  937] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  938] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  939] = 32'b11000010110111100000000000000000;
	assign	noise_gru_recurrent_weights_array[  940] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  941] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  942] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  943] = 32'b11000010110001100000000000000000;
	assign	noise_gru_recurrent_weights_array[  944] = 32'b11000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[  945] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  946] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  947] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  948] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  949] = 32'b11000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  950] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  951] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  952] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  953] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  954] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  955] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  956] = 32'b01000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  957] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  958] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  959] = 32'b01000010110111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  960] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  961] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  962] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  963] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[  964] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  965] = 32'b11000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[  966] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  967] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  968] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  969] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  970] = 32'b11000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[  971] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  972] = 32'b11000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[  973] = 32'b11000011000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  974] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  975] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  976] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  977] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  978] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  979] = 32'b01000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  980] = 32'b11000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[  981] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[  982] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  983] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  984] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  985] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[  986] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  987] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  988] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  989] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  990] = 32'b11000010110101100000000000000000;
	assign	noise_gru_recurrent_weights_array[  991] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  992] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[  993] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  994] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[  995] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[  996] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[  997] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[  998] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[  999] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1000] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1001] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1002] = 32'b11000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1003] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1004] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1005] = 32'b01000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1006] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1007] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1008] = 32'b11000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1009] = 32'b11000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1010] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1011] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1012] = 32'b11000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1013] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1014] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1015] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1016] = 32'b11000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1017] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1018] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1019] = 32'b01000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1020] = 32'b11000010110111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1021] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1022] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1023] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1024] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1025] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1026] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1027] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1028] = 32'b01000010110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1029] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1030] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1031] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1032] = 32'b01000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1033] = 32'b11000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1034] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1035] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1036] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1037] = 32'b01000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1038] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1039] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1040] = 32'b11000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1041] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1042] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1043] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1044] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1045] = 32'b01000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1046] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1047] = 32'b11000010110111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1048] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1049] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1050] = 32'b01000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1051] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1052] = 32'b01000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1053] = 32'b01000010110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1054] = 32'b11000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1055] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1056] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1057] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1058] = 32'b01000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1059] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1060] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1061] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1062] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1063] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1064] = 32'b11000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1065] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1066] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1067] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1068] = 32'b01000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1069] = 32'b11000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1070] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1071] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1072] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1073] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1074] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1075] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1076] = 32'b11000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1077] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1078] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1079] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1080] = 32'b01000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1081] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1082] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1083] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1084] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1085] = 32'b01000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1086] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1087] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1088] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1089] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1090] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1091] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1092] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1093] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1094] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1095] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1096] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1097] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1098] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1099] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1100] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1101] = 32'b01000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1102] = 32'b11000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1103] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1104] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1105] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1106] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1107] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1108] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1109] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1110] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1111] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1112] = 32'b01000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1113] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1114] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1115] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1116] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1117] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1118] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1119] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1120] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1121] = 32'b11000010110100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1122] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1123] = 32'b01000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1124] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1125] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1126] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1127] = 32'b01000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1128] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1129] = 32'b11000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1130] = 32'b01000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1131] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1132] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1133] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1134] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1135] = 32'b01000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1136] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1137] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1138] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1139] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1140] = 32'b01000010110100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1141] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1142] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1143] = 32'b11000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1144] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1145] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1146] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1147] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1148] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1149] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1150] = 32'b01000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1151] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1152] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1153] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1154] = 32'b01000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1155] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1156] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1157] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1158] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1159] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1160] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1161] = 32'b01000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1162] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1163] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1164] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1165] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1166] = 32'b11000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1167] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1168] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1169] = 32'b01000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1170] = 32'b11000010110111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1171] = 32'b11000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1172] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1173] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1174] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1175] = 32'b01000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1176] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1177] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1178] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1179] = 32'b01000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1180] = 32'b01000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1181] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1182] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1183] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1184] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1185] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1186] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1187] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1188] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1189] = 32'b11000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1190] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1191] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1192] = 32'b01000010101100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1193] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1194] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1195] = 32'b01000010111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1196] = 32'b11000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1197] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1198] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1199] = 32'b01000010111001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1200] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1201] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1202] = 32'b11000010110011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1203] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1204] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1205] = 32'b01000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1206] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1207] = 32'b11000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1208] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1209] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1210] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1211] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1212] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1213] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1214] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1215] = 32'b11000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1216] = 32'b01000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1217] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1218] = 32'b11000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1219] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1220] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1221] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1222] = 32'b01000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1223] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1224] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1225] = 32'b01000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1226] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1227] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1228] = 32'b01000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1229] = 32'b01000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1230] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1231] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1232] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1233] = 32'b01000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1234] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1235] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1236] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1237] = 32'b11000010110101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1238] = 32'b01000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1239] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1240] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1241] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1242] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1243] = 32'b11000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1244] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1245] = 32'b11000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1246] = 32'b01000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1247] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1248] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1249] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1250] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1251] = 32'b01000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1252] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1253] = 32'b01000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1254] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1255] = 32'b01000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1256] = 32'b01000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1257] = 32'b01000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1258] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1259] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1260] = 32'b11000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1261] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1262] = 32'b11000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1263] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1264] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1265] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1266] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1267] = 32'b11000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1268] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1269] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1270] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1271] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1272] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1273] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1274] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1275] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1276] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1277] = 32'b01000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1278] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1279] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1280] = 32'b11000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1281] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1282] = 32'b11000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1283] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1284] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1285] = 32'b01000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1286] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1287] = 32'b11000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1288] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1289] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1290] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1291] = 32'b01000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1292] = 32'b01000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1293] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1294] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1295] = 32'b01000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1296] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1297] = 32'b11000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1298] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1299] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1300] = 32'b11000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1301] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1302] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1303] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1304] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1305] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1306] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1307] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1308] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1309] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1310] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1311] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1312] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1313] = 32'b11000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1314] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1315] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1316] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1317] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1318] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1319] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1320] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1321] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1322] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1323] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1324] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1325] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1326] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1327] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1328] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1329] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1330] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1331] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1332] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1333] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1334] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1335] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1336] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1337] = 32'b11000010111001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1338] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1339] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1340] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1341] = 32'b01000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1342] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1343] = 32'b01000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1344] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1345] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1346] = 32'b01000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1347] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1348] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1349] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1350] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1351] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1352] = 32'b11000010110111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1353] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1354] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1355] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1356] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1357] = 32'b11000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1358] = 32'b11000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1359] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1360] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1361] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1362] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1363] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1364] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1365] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1366] = 32'b01000010110101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1367] = 32'b01000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1368] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1369] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1370] = 32'b01000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1371] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1372] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1373] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1374] = 32'b01000010110011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1375] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1376] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1377] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1378] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1379] = 32'b11000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1380] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1381] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1382] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1383] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1384] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1385] = 32'b01000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1386] = 32'b11000010110101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1387] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1388] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1389] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1390] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1391] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1392] = 32'b11000010110111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1393] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1394] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1395] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1396] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1397] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1398] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1399] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1400] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1401] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1402] = 32'b11000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1403] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1404] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1405] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1406] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1407] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1408] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1409] = 32'b01000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1410] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1411] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1412] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1413] = 32'b11000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1414] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1415] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1416] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1417] = 32'b11000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1418] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1419] = 32'b01000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1420] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1421] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1422] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1423] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1424] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1425] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1426] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1427] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1428] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1429] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1430] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1431] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1432] = 32'b11000010110101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1433] = 32'b01000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1434] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1435] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1436] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1437] = 32'b11000010110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1438] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1439] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1440] = 32'b11000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1441] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1442] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1443] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1444] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1445] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1446] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1447] = 32'b11000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1448] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1449] = 32'b01000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1450] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1451] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1452] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1453] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1454] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1455] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1456] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1457] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1458] = 32'b01000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1459] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1460] = 32'b01000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1461] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1462] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1463] = 32'b01000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1464] = 32'b01000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1465] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1466] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1467] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1468] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1469] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1470] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1471] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1472] = 32'b11000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1473] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1474] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1475] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1476] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1477] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1478] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1479] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1480] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1481] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1482] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1483] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1484] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1485] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1486] = 32'b11000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1487] = 32'b11000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1488] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1489] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1490] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1491] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1492] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1493] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1494] = 32'b01000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1495] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1496] = 32'b11000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1497] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1498] = 32'b11000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1499] = 32'b01000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1500] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1501] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1502] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1503] = 32'b01000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1504] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1505] = 32'b01000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1506] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1507] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1508] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1509] = 32'b01000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1510] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1511] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1512] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1513] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1514] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1515] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1516] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1517] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1518] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1519] = 32'b11000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1520] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1521] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1522] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1523] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1524] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1525] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1526] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1527] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1528] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1529] = 32'b11000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1530] = 32'b01000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1531] = 32'b11000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1532] = 32'b11000010111001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1533] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1534] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1535] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1536] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1537] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1538] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1539] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1540] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1541] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1542] = 32'b11000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1543] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1544] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1545] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1546] = 32'b01000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1547] = 32'b11000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1548] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1549] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1550] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1551] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1552] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1553] = 32'b11000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1554] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1555] = 32'b01000010101110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1556] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1557] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1558] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1559] = 32'b11000011000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1560] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1561] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1562] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1563] = 32'b11000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1564] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1565] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1566] = 32'b11000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1567] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1568] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1569] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1570] = 32'b01000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1571] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1572] = 32'b11000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1573] = 32'b11000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1574] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1575] = 32'b01000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1576] = 32'b01000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1577] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1578] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1579] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1580] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1581] = 32'b11000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1582] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1583] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1584] = 32'b11000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1585] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1586] = 32'b11000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1587] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1588] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1589] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1590] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1591] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1592] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1593] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1594] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1595] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1596] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1597] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1598] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1599] = 32'b11000010110011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1600] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1601] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1602] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1603] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1604] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1605] = 32'b01000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1606] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1607] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1608] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1609] = 32'b11000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1610] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1611] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1612] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1613] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1614] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1615] = 32'b11000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1616] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1617] = 32'b01000010110001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1618] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1619] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1620] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1621] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1622] = 32'b01000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1623] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1624] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1625] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1626] = 32'b11000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1627] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1628] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1629] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1630] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1631] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1632] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1633] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1634] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1635] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1636] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1637] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1638] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1639] = 32'b11000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1640] = 32'b11000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1641] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1642] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1643] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1644] = 32'b01000010110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1645] = 32'b01000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1646] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1647] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1648] = 32'b01000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1649] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1650] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1651] = 32'b01000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1652] = 32'b01000010111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1653] = 32'b11000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1654] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1655] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1656] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1657] = 32'b11000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1658] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1659] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1660] = 32'b01000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1661] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1662] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1663] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1664] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1665] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1666] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1667] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1668] = 32'b01000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1669] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1670] = 32'b01000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1671] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1672] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1673] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1674] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1675] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1676] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1677] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1678] = 32'b01000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1679] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1680] = 32'b11000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1681] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1682] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1683] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1684] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1685] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1686] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1687] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1688] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1689] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1690] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1691] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1692] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1693] = 32'b01000010110100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1694] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1695] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1696] = 32'b01000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1697] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1698] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1699] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1700] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1701] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1702] = 32'b01000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1703] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1704] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1705] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1706] = 32'b01000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1707] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1708] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1709] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1710] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1711] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1712] = 32'b11000010101110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1713] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1714] = 32'b11000010110101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1715] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1716] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1717] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1718] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1719] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1720] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1721] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1722] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1723] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1724] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1725] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1726] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1727] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1728] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1729] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1730] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1731] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1732] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1733] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1734] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1735] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1736] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1737] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1738] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1739] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1740] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1741] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1742] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1743] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1744] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1745] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1746] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1747] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1748] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1749] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1750] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1751] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1752] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1753] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1754] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1755] = 32'b01000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1756] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1757] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1758] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1759] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1760] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1761] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1762] = 32'b01000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1763] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1764] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1765] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1766] = 32'b01000010111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1767] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1768] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1769] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1770] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1771] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1772] = 32'b01000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1773] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1774] = 32'b01000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1775] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1776] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1777] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1778] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1779] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1780] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1781] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1782] = 32'b01000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1783] = 32'b11000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1784] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1785] = 32'b11000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1786] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1787] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1788] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1789] = 32'b11000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1790] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1791] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1792] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1793] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1794] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1795] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1796] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1797] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1798] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1799] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1800] = 32'b01000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1801] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1802] = 32'b11000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1803] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1804] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1805] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1806] = 32'b01000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1807] = 32'b11000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1808] = 32'b01000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1809] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1810] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1811] = 32'b11000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1812] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1813] = 32'b11000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1814] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1815] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1816] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1817] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1818] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1819] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1820] = 32'b01000010110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1821] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1822] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1823] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1824] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1825] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1826] = 32'b11000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1827] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1828] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1829] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1830] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1831] = 32'b01000010110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1832] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1833] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1834] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1835] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1836] = 32'b11000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1837] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1838] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1839] = 32'b01000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1840] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1841] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1842] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1843] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1844] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1845] = 32'b01000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1846] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1847] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1848] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1849] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1850] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1851] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1852] = 32'b11000010111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1853] = 32'b11000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1854] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1855] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1856] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1857] = 32'b11000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1858] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1859] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1860] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1861] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1862] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1863] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1864] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1865] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1866] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1867] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1868] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1869] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1870] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1871] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1872] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1873] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1874] = 32'b01000010110111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1875] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1876] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1877] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1878] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1879] = 32'b01000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1880] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1881] = 32'b01000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1882] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1883] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1884] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1885] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1886] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1887] = 32'b01000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1888] = 32'b01000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1889] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1890] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1891] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1892] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1893] = 32'b11000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1894] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1895] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1896] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1897] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1898] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1899] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1900] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1901] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1902] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1903] = 32'b01000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1904] = 32'b01000010110111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1905] = 32'b11000010110100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1906] = 32'b01000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1907] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1908] = 32'b01000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1909] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1910] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1911] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1912] = 32'b01000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1913] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1914] = 32'b01000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1915] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1916] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1917] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1918] = 32'b01000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1919] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1920] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1921] = 32'b11000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1922] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1923] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1924] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1925] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1926] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1927] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1928] = 32'b11000010110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1929] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1930] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1931] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1932] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1933] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1934] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1935] = 32'b11000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1936] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1937] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1938] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1939] = 32'b11000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1940] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1941] = 32'b01000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1942] = 32'b11000010110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1943] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1944] = 32'b01000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1945] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1946] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1947] = 32'b01000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1948] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1949] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1950] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1951] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1952] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1953] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1954] = 32'b11000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1955] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1956] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1957] = 32'b01000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1958] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1959] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1960] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1961] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1962] = 32'b01000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1963] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1964] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1965] = 32'b01000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1966] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1967] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1968] = 32'b01000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1969] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1970] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1971] = 32'b01000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1972] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1973] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1974] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1975] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1976] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1977] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1978] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1979] = 32'b01000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1980] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1981] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1982] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1983] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1984] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1985] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1986] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1987] = 32'b01000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1988] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1989] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1990] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1991] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1992] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1993] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1994] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1995] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1996] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1997] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1998] = 32'b11000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 1999] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2000] = 32'b11000010110001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2001] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2002] = 32'b01000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2003] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2004] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2005] = 32'b11000010110011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2006] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2007] = 32'b11000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2008] = 32'b11000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2009] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2010] = 32'b01000010110001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2011] = 32'b11000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2012] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2013] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2014] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2015] = 32'b11000010110111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2016] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2017] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2018] = 32'b11000010110001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2019] = 32'b11000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2020] = 32'b01000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2021] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2022] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2023] = 32'b01000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2024] = 32'b11000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2025] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2026] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2027] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2028] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2029] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2030] = 32'b11000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2031] = 32'b11000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2032] = 32'b01000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2033] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2034] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2035] = 32'b01000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2036] = 32'b11000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2037] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2038] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2039] = 32'b11000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2040] = 32'b11000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2041] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2042] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2043] = 32'b11000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2044] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2045] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2046] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2047] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2048] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2049] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2050] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2051] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2052] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2053] = 32'b01000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2054] = 32'b11000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2055] = 32'b01000010111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2056] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2057] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2058] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2059] = 32'b01000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2060] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2061] = 32'b11000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2062] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2063] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2064] = 32'b11000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2065] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2066] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2067] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2068] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2069] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2070] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2071] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2072] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2073] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2074] = 32'b11000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2075] = 32'b01000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2076] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2077] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2078] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2079] = 32'b01000010110001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2080] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2081] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2082] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2083] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2084] = 32'b11000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2085] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2086] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2087] = 32'b11000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2088] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2089] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2090] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2091] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2092] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2093] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2094] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2095] = 32'b11000010110111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2096] = 32'b01000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2097] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2098] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2099] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2100] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2101] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2102] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2103] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2104] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2105] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2106] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2107] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2108] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2109] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2110] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2111] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2112] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2113] = 32'b01000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2114] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2115] = 32'b01000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2116] = 32'b11000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2117] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2118] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2119] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2120] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2121] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2122] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2123] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2124] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2125] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2126] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2127] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2128] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2129] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2130] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2131] = 32'b01000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2132] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2133] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2134] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2135] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2136] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2137] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2138] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2139] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2140] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2141] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2142] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2143] = 32'b11000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2144] = 32'b11000010110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2145] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2146] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2147] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2148] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2149] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2150] = 32'b11000010110111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2151] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2152] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2153] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2154] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2155] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2156] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2157] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2158] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2159] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2160] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2161] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2162] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2163] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2164] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2165] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2166] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2167] = 32'b01000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2168] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2169] = 32'b01000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2170] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2171] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2172] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2173] = 32'b01000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2174] = 32'b01000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2175] = 32'b01000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2176] = 32'b01000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2177] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2178] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2179] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2180] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2181] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2182] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2183] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2184] = 32'b01000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2185] = 32'b01000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2186] = 32'b01000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2187] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2188] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2189] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2190] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2191] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2192] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2193] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2194] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2195] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2196] = 32'b11000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2197] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2198] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2199] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2200] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2201] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2202] = 32'b01000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2203] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2204] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2205] = 32'b01000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2206] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2207] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2208] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2209] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2210] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2211] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2212] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2213] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2214] = 32'b11000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2215] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2216] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2217] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2218] = 32'b11000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2219] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2220] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2221] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2222] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2223] = 32'b01000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2224] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2225] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2226] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2227] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2228] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2229] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2230] = 32'b01000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2231] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2232] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2233] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2234] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2235] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2236] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2237] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2238] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2239] = 32'b01000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2240] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2241] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2242] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2243] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2244] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2245] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2246] = 32'b01000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2247] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2248] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2249] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2250] = 32'b01000010110101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2251] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2252] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2253] = 32'b01000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2254] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2255] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2256] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2257] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2258] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2259] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2260] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2261] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2262] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2263] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2264] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2265] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2266] = 32'b01000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2267] = 32'b01000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2268] = 32'b11000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2269] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2270] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2271] = 32'b11000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2272] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2273] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2274] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2275] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2276] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2277] = 32'b11000010110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2278] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2279] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2280] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2281] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2282] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2283] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2284] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2285] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2286] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2287] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2288] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2289] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2290] = 32'b01000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2291] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2292] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2293] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2294] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2295] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2296] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2297] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2298] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2299] = 32'b01000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2300] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2301] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2302] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2303] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2304] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2305] = 32'b11000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2306] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2307] = 32'b01000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2308] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2309] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2310] = 32'b11000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2311] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2312] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2313] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2314] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2315] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2316] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2317] = 32'b01000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2318] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2319] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2320] = 32'b01000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2321] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2322] = 32'b01000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2323] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2324] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2325] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2326] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2327] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2328] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2329] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2330] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2331] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2332] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2333] = 32'b01000010110111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2334] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2335] = 32'b11000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2336] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2337] = 32'b01000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2338] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2339] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2340] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2341] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2342] = 32'b01000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2343] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2344] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2345] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2346] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2347] = 32'b11000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2348] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2349] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2350] = 32'b01000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2351] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2352] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2353] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2354] = 32'b01000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2355] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2356] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2357] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2358] = 32'b01000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2359] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2360] = 32'b11000010110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2361] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2362] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2363] = 32'b11000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2364] = 32'b01000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2365] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2366] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2367] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2368] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2369] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2370] = 32'b11000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2371] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2372] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2373] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2374] = 32'b11000010110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2375] = 32'b11000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2376] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2377] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2378] = 32'b01000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2379] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2380] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2381] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2382] = 32'b01000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2383] = 32'b11000010110101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2384] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2385] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2386] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2387] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2388] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2389] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2390] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2391] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2392] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2393] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2394] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2395] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2396] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2397] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2398] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2399] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2400] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2401] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2402] = 32'b11000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2403] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2404] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2405] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2406] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2407] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2408] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2409] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2410] = 32'b11000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2411] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2412] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2413] = 32'b01000010111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2414] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2415] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2416] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2417] = 32'b11000010111001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2418] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2419] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2420] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2421] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2422] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2423] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2424] = 32'b01000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2425] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2426] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2427] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2428] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2429] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2430] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2431] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2432] = 32'b11000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2433] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2434] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2435] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2436] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2437] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2438] = 32'b01000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2439] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2440] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2441] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2442] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2443] = 32'b11000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2444] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2445] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2446] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2447] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2448] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2449] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2450] = 32'b01000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2451] = 32'b01000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2452] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2453] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2454] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2455] = 32'b01000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2456] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2457] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2458] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2459] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2460] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2461] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2462] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2463] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2464] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2465] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2466] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2467] = 32'b01000010110100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2468] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2469] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2470] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2471] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2472] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2473] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2474] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2475] = 32'b01000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2476] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2477] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2478] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2479] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2480] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2481] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2482] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2483] = 32'b01000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2484] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2485] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2486] = 32'b01000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2487] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2488] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2489] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2490] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2491] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2492] = 32'b11000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2493] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2494] = 32'b01000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2495] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2496] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2497] = 32'b01000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2498] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2499] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2500] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2501] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2502] = 32'b01000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2503] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2504] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2505] = 32'b11000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2506] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2507] = 32'b11000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2508] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2509] = 32'b01000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2510] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2511] = 32'b01000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2512] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2513] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2514] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2515] = 32'b01000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2516] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2517] = 32'b11000010110001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2518] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2519] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2520] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2521] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2522] = 32'b01000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2523] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2524] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2525] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2526] = 32'b11000011000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2527] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2528] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2529] = 32'b11000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2530] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2531] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2532] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2533] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2534] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2535] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2536] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2537] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2538] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2539] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2540] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2541] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2542] = 32'b11000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2543] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2544] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2545] = 32'b11000010101110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2546] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2547] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2548] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2549] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2550] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2551] = 32'b11000010110111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2552] = 32'b01000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2553] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2554] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2555] = 32'b11000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2556] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2557] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2558] = 32'b01000010110101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2559] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2560] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2561] = 32'b01000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2562] = 32'b11000010110011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2563] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2564] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2565] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2566] = 32'b11000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2567] = 32'b01000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2568] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2569] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2570] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2571] = 32'b11000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2572] = 32'b01000010110101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2573] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2574] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2575] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2576] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2577] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2578] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2579] = 32'b11000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2580] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2581] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2582] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2583] = 32'b11000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2584] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2585] = 32'b01000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2586] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2587] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2588] = 32'b11000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2589] = 32'b01000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2590] = 32'b11000010111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2591] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2592] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2593] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2594] = 32'b01000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2595] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2596] = 32'b11000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2597] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2598] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2599] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2600] = 32'b11000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2601] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2602] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2603] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2604] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2605] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2606] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2607] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2608] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2609] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2610] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2611] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2612] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2613] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2614] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2615] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2616] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2617] = 32'b11000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2618] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2619] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2620] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2621] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2622] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2623] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2624] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2625] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2626] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2627] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2628] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2629] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2630] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2631] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2632] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2633] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2634] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2635] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2636] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2637] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2638] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2639] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2640] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2641] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2642] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2643] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2644] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2645] = 32'b01000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2646] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2647] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2648] = 32'b01000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2649] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2650] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2651] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2652] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2653] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2654] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2655] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2656] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2657] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2658] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2659] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2660] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2661] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2662] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2663] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2664] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2665] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2666] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2667] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2668] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2669] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2670] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2671] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2672] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2673] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2674] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2675] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2676] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2677] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2678] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2679] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2680] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2681] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2682] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2683] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2684] = 32'b11000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2685] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2686] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2687] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2688] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2689] = 32'b01000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2690] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2691] = 32'b01000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2692] = 32'b11000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2693] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2694] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2695] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2696] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2697] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2698] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2699] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2700] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2701] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2702] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2703] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2704] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2705] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2706] = 32'b11000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2707] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2708] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2709] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2710] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2711] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2712] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2713] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2714] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2715] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2716] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2717] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2718] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2719] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2720] = 32'b01000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2721] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2722] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2723] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2724] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2725] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2726] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2727] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2728] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2729] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2730] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2731] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2732] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2733] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2734] = 32'b01000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2735] = 32'b11000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2736] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2737] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2738] = 32'b01000010110011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2739] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2740] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2741] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2742] = 32'b11000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2743] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2744] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2745] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2746] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2747] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2748] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2749] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2750] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2751] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2752] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2753] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2754] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2755] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2756] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2757] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2758] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2759] = 32'b01000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2760] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2761] = 32'b11000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2762] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2763] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2764] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2765] = 32'b11000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2766] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2767] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2768] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2769] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2770] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2771] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2772] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2773] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2774] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2775] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2776] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2777] = 32'b11000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2778] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2779] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2780] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2781] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2782] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2783] = 32'b01000010110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2784] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2785] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2786] = 32'b01000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2787] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2788] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2789] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2790] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2791] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2792] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2793] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2794] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2795] = 32'b01000010110111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2796] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2797] = 32'b11000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2798] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2799] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2800] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2801] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2802] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2803] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2804] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2805] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2806] = 32'b11000010101110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2807] = 32'b01000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2808] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2809] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2810] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2811] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2812] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2813] = 32'b11000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2814] = 32'b01000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2815] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2816] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2817] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2818] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2819] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2820] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2821] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2822] = 32'b11000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2823] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2824] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2825] = 32'b11000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2826] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2827] = 32'b11000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2828] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2829] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2830] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2831] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2832] = 32'b01000010110101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2833] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2834] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2835] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2836] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2837] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2838] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2839] = 32'b01000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2840] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2841] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2842] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2843] = 32'b11000010101100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2844] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2845] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2846] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2847] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2848] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2849] = 32'b11000010111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2850] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2851] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2852] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2853] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2854] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2855] = 32'b11000010111001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2856] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2857] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2858] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2859] = 32'b11000010110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2860] = 32'b11000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2861] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2862] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2863] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2864] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2865] = 32'b11000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2866] = 32'b11000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2867] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2868] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2869] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2870] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2871] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2872] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2873] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2874] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2875] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2876] = 32'b11000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2877] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2878] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2879] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2880] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2881] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2882] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2883] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2884] = 32'b01000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2885] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2886] = 32'b11000010110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2887] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2888] = 32'b01000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2889] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2890] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2891] = 32'b01000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2892] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2893] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2894] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2895] = 32'b01000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2896] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2897] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2898] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2899] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2900] = 32'b11000011000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2901] = 32'b01000010110111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2902] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2903] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2904] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2905] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2906] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2907] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2908] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2909] = 32'b01000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2910] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2911] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2912] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2913] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2914] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2915] = 32'b01000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2916] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2917] = 32'b01000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2918] = 32'b01000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2919] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2920] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2921] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2922] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2923] = 32'b11000010110001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2924] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2925] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2926] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2927] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2928] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2929] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2930] = 32'b11000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2931] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2932] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2933] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2934] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2935] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2936] = 32'b11000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2937] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2938] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2939] = 32'b01000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2940] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2941] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2942] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2943] = 32'b01000010110111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2944] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2945] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2946] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2947] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2948] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2949] = 32'b01000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2950] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2951] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2952] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2953] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2954] = 32'b01000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2955] = 32'b01000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2956] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2957] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2958] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2959] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2960] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2961] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2962] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2963] = 32'b11000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2964] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2965] = 32'b01000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2966] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2967] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2968] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2969] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2970] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2971] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2972] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2973] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2974] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2975] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2976] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2977] = 32'b01000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2978] = 32'b11000010110011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2979] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2980] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2981] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2982] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2983] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2984] = 32'b11000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2985] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2986] = 32'b11000011000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2987] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2988] = 32'b11000010110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2989] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2990] = 32'b01000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2991] = 32'b01000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2992] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2993] = 32'b11000011000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2994] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2995] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2996] = 32'b11000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2997] = 32'b11000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2998] = 32'b01000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 2999] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3000] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3001] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3002] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3003] = 32'b11000010101110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3004] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3005] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3006] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3007] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3008] = 32'b11000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3009] = 32'b11000010110111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3010] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3011] = 32'b11000010110100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3012] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3013] = 32'b11000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3014] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3015] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3016] = 32'b11000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3017] = 32'b11000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3018] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3019] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3020] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3021] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3022] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3023] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3024] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3025] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3026] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3027] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3028] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3029] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3030] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3031] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3032] = 32'b11000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3033] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3034] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3035] = 32'b01000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3036] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3037] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3038] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3039] = 32'b01000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3040] = 32'b01000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3041] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3042] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3043] = 32'b01000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3044] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3045] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3046] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3047] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3048] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3049] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3050] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3051] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3052] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3053] = 32'b01000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3054] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3055] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3056] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3057] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3058] = 32'b01000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3059] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3060] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3061] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3062] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3063] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3064] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3065] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3066] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3067] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3068] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3069] = 32'b01000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3070] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3071] = 32'b01000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3072] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3073] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3074] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3075] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3076] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3077] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3078] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3079] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3080] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3081] = 32'b01000010110011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3082] = 32'b11000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3083] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3084] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3085] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3086] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3087] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3088] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3089] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3090] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3091] = 32'b11000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3092] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3093] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3094] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3095] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3096] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3097] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3098] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3099] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3100] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3101] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3102] = 32'b11000010111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3103] = 32'b11000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3104] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3105] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3106] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3107] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3108] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3109] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3110] = 32'b01000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3111] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3112] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3113] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3114] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3115] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3116] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3117] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3118] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3119] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3120] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3121] = 32'b11000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3122] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3123] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3124] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3125] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3126] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3127] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3128] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3129] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3130] = 32'b11000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3131] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3132] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3133] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3134] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3135] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3136] = 32'b01000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3137] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3138] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3139] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3140] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3141] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3142] = 32'b11000010111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3143] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3144] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3145] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3146] = 32'b01000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3147] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3148] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3149] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3150] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3151] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3152] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3153] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3154] = 32'b11000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3155] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3156] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3157] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3158] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3159] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3160] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3161] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3162] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3163] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3164] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3165] = 32'b11000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3166] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3167] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3168] = 32'b11000010110001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3169] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3170] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3171] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3172] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3173] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3174] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3175] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3176] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3177] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3178] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3179] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3180] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3181] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3182] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3183] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3184] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3185] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3186] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3187] = 32'b11000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3188] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3189] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3190] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3191] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3192] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3193] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3194] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3195] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3196] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3197] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3198] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3199] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3200] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3201] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3202] = 32'b01000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3203] = 32'b11000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3204] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3205] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3206] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3207] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3208] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3209] = 32'b01000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3210] = 32'b01000010110100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3211] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3212] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3213] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3214] = 32'b01000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3215] = 32'b01000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3216] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3217] = 32'b11000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3218] = 32'b11000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3219] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3220] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3221] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3222] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3223] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3224] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3225] = 32'b01000010110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3226] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3227] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3228] = 32'b11000010101100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3229] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3230] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3231] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3232] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3233] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3234] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3235] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3236] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3237] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3238] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3239] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3240] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3241] = 32'b01000010101100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3242] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3243] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3244] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3245] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3246] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3247] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3248] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3249] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3250] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3251] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3252] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3253] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3254] = 32'b11000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3255] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3256] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3257] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3258] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3259] = 32'b01000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3260] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3261] = 32'b11000010111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3262] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3263] = 32'b11000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3264] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3265] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3266] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3267] = 32'b01000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3268] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3269] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3270] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3271] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3272] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3273] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3274] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3275] = 32'b11000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3276] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3277] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3278] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3279] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3280] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3281] = 32'b01000010110111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3282] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3283] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3284] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3285] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3286] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3287] = 32'b11000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3288] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3289] = 32'b01000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3290] = 32'b11000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3291] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3292] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3293] = 32'b01000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3294] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3295] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3296] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3297] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3298] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3299] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3300] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3301] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3302] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3303] = 32'b11000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3304] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3305] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3306] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3307] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3308] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3309] = 32'b11000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3310] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3311] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3312] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3313] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3314] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3315] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3316] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3317] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3318] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3319] = 32'b01000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3320] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3321] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3322] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3323] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3324] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3325] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3326] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3327] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3328] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3329] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3330] = 32'b01000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3331] = 32'b01000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3332] = 32'b01000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3333] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3334] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3335] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3336] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3337] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3338] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3339] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3340] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3341] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3342] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3343] = 32'b11000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3344] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3345] = 32'b01000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3346] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3347] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3348] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3349] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3350] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3351] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3352] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3353] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3354] = 32'b01000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3355] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3356] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3357] = 32'b01000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3358] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3359] = 32'b01000010110011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3360] = 32'b11000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3361] = 32'b01000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3362] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3363] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3364] = 32'b01000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3365] = 32'b01000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3366] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3367] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3368] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3369] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3370] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3371] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3372] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3373] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3374] = 32'b01000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3375] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3376] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3377] = 32'b01000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3378] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3379] = 32'b11000010110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3380] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3381] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3382] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3383] = 32'b11000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3384] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3385] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3386] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3387] = 32'b01000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3388] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3389] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3390] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3391] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3392] = 32'b01000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3393] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3394] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3395] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3396] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3397] = 32'b11000011000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3398] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3399] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3400] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3401] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3402] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3403] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3404] = 32'b01000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3405] = 32'b11000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3406] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3407] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3408] = 32'b11000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3409] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3410] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3411] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3412] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3413] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3414] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3415] = 32'b01000010110111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3416] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3417] = 32'b01000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3418] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3419] = 32'b11000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3420] = 32'b01000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3421] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3422] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3423] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3424] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3425] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3426] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3427] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3428] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3429] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3430] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3431] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3432] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3433] = 32'b11000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3434] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3435] = 32'b11000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3436] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3437] = 32'b01000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3438] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3439] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3440] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3441] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3442] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3443] = 32'b11000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3444] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3445] = 32'b01000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3446] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3447] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3448] = 32'b01000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3449] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3450] = 32'b01000010101100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3451] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3452] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3453] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3454] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3455] = 32'b01000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3456] = 32'b11000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3457] = 32'b11000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3458] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3459] = 32'b11000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3460] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3461] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3462] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3463] = 32'b01000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3464] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3465] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3466] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3467] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3468] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3469] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3470] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3471] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3472] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3473] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3474] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3475] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3476] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3477] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3478] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3479] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3480] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3481] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3482] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3483] = 32'b01000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3484] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3485] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3486] = 32'b01000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3487] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3488] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3489] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3490] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3491] = 32'b01000010110100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3492] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3493] = 32'b11000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3494] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3495] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3496] = 32'b01000010110011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3497] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3498] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3499] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3500] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3501] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3502] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3503] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3504] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3505] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3506] = 32'b01000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3507] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3508] = 32'b01000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3509] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3510] = 32'b01000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3511] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3512] = 32'b01000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3513] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3514] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3515] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3516] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3517] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3518] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3519] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3520] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3521] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3522] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3523] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3524] = 32'b11000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3525] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3526] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3527] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3528] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3529] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3530] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3531] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3532] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3533] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3534] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3535] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3536] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3537] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3538] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3539] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3540] = 32'b01000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3541] = 32'b11000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3542] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3543] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3544] = 32'b11000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3545] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3546] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3547] = 32'b11000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3548] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3549] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3550] = 32'b11000010110111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3551] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3552] = 32'b01000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3553] = 32'b01000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3554] = 32'b01000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3555] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3556] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3557] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3558] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3559] = 32'b11000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3560] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3561] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3562] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3563] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3564] = 32'b11000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3565] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3566] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3567] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3568] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3569] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3570] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3571] = 32'b01000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3572] = 32'b01000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3573] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3574] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3575] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3576] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3577] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3578] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3579] = 32'b01000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3580] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3581] = 32'b01000010110101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3582] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3583] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3584] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3585] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3586] = 32'b01000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3587] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3588] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3589] = 32'b11000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3590] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3591] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3592] = 32'b11000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3593] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3594] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3595] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3596] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3597] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3598] = 32'b11000011000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3599] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3600] = 32'b11000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3601] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3602] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3603] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3604] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3605] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3606] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3607] = 32'b01000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3608] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3609] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3610] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3611] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3612] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3613] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3614] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3615] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3616] = 32'b01000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3617] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3618] = 32'b01000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3619] = 32'b01000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3620] = 32'b11000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3621] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3622] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3623] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3624] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3625] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3626] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3627] = 32'b01000010110001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3628] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3629] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3630] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3631] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3632] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3633] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3634] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3635] = 32'b01000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3636] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3637] = 32'b01000010110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3638] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3639] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3640] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3641] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3642] = 32'b11000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3643] = 32'b11000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3644] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3645] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3646] = 32'b01000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3647] = 32'b11000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3648] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3649] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3650] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3651] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3652] = 32'b01000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3653] = 32'b01000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3654] = 32'b01000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3655] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3656] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3657] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3658] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3659] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3660] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3661] = 32'b01000010101100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3662] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3663] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3664] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3665] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3666] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3667] = 32'b11000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3668] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3669] = 32'b11000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3670] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3671] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3672] = 32'b01000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3673] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3674] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3675] = 32'b01000010110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3676] = 32'b11000010110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3677] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3678] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3679] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3680] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3681] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3682] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3683] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3684] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3685] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3686] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3687] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3688] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3689] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3690] = 32'b11000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3691] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3692] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3693] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3694] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3695] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3696] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3697] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3698] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3699] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3700] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3701] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3702] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3703] = 32'b11000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3704] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3705] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3706] = 32'b01000010110101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3707] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3708] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3709] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3710] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3711] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3712] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3713] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3714] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3715] = 32'b11000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3716] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3717] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3718] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3719] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3720] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3721] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3722] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3723] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3724] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3725] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3726] = 32'b01000010101100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3727] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3728] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3729] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3730] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3731] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3732] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3733] = 32'b11000011000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3734] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3735] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3736] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3737] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3738] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3739] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3740] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3741] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3742] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3743] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3744] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3745] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3746] = 32'b01000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3747] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3748] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3749] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3750] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3751] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3752] = 32'b01000010110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3753] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3754] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3755] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3756] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3757] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3758] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3759] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3760] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3761] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3762] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3763] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3764] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3765] = 32'b01000010110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3766] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3767] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3768] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3769] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3770] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3771] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3772] = 32'b01000010110001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3773] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3774] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3775] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3776] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3777] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3778] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3779] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3780] = 32'b01000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3781] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3782] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3783] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3784] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3785] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3786] = 32'b01000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3787] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3788] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3789] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3790] = 32'b01000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3791] = 32'b01000010110001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3792] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3793] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3794] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3795] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3796] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3797] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3798] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3799] = 32'b11000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3800] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3801] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3802] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3803] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3804] = 32'b01000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3805] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3806] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3807] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3808] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3809] = 32'b01000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3810] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3811] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3812] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3813] = 32'b01000010110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3814] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3815] = 32'b11000010110101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3816] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3817] = 32'b01000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3818] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3819] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3820] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3821] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3822] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3823] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3824] = 32'b11000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3825] = 32'b01000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3826] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3827] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3828] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3829] = 32'b11000010111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3830] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3831] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3832] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3833] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3834] = 32'b11000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3835] = 32'b01000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3836] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3837] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3838] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3839] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3840] = 32'b01000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3841] = 32'b11000010110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3842] = 32'b01000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3843] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3844] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3845] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3846] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3847] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3848] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3849] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3850] = 32'b11000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3851] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3852] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3853] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3854] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3855] = 32'b01000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3856] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3857] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3858] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3859] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3860] = 32'b11000010101110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3861] = 32'b11000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3862] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3863] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3864] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3865] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3866] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3867] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3868] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3869] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3870] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3871] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3872] = 32'b11000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3873] = 32'b01000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3874] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3875] = 32'b11000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3876] = 32'b11000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3877] = 32'b11000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3878] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3879] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3880] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3881] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3882] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3883] = 32'b11000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3884] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3885] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3886] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3887] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3888] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3889] = 32'b01000010110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3890] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3891] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3892] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3893] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3894] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3895] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3896] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3897] = 32'b01000010110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3898] = 32'b01000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3899] = 32'b01000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3900] = 32'b01000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3901] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3902] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3903] = 32'b01000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3904] = 32'b01000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3905] = 32'b11000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3906] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3907] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3908] = 32'b01000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3909] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3910] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3911] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3912] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3913] = 32'b01000010110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3914] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3915] = 32'b01000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3916] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3917] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3918] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3919] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3920] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3921] = 32'b01000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3922] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3923] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3924] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3925] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3926] = 32'b01000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3927] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3928] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3929] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3930] = 32'b01000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3931] = 32'b11000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3932] = 32'b01000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3933] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3934] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3935] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3936] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3937] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3938] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3939] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3940] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3941] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3942] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3943] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3944] = 32'b01000010111001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3945] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3946] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3947] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3948] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3949] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3950] = 32'b01000010110111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3951] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3952] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3953] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3954] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3955] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3956] = 32'b01000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3957] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3958] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3959] = 32'b01000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3960] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3961] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3962] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3963] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3964] = 32'b01000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3965] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3966] = 32'b11000010110011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3967] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3968] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3969] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3970] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3971] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3972] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3973] = 32'b01000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3974] = 32'b01000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3975] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3976] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3977] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3978] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3979] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3980] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3981] = 32'b11000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3982] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3983] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3984] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3985] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3986] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3987] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3988] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3989] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3990] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3991] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3992] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3993] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3994] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3995] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3996] = 32'b01000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3997] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3998] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 3999] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4000] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4001] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4002] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4003] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4004] = 32'b11000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4005] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4006] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4007] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4008] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4009] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4010] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4011] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4012] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4013] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4014] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4015] = 32'b01000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4016] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4017] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4018] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4019] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4020] = 32'b11000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4021] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4022] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4023] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4024] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4025] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4026] = 32'b11000010110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4027] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4028] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4029] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4030] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4031] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4032] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4033] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4034] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4035] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4036] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4037] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4038] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4039] = 32'b01000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4040] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4041] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4042] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4043] = 32'b01000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4044] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4045] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4046] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4047] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4048] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4049] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4050] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4051] = 32'b11000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4052] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4053] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4054] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4055] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4056] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4057] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4058] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4059] = 32'b01000010110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4060] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4061] = 32'b01000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4062] = 32'b01000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4063] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4064] = 32'b11000010110100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4065] = 32'b11000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4066] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4067] = 32'b01000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4068] = 32'b11000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4069] = 32'b01000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4070] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4071] = 32'b11000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4072] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4073] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4074] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4075] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4076] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4077] = 32'b11000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4078] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4079] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4080] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4081] = 32'b11000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4082] = 32'b01000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4083] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4084] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4085] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4086] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4087] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4088] = 32'b01000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4089] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4090] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4091] = 32'b11000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4092] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4093] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4094] = 32'b01000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4095] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4096] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4097] = 32'b01000010110111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4098] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4099] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4100] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4101] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4102] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4103] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4104] = 32'b01000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4105] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4106] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4107] = 32'b11000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4108] = 32'b11000010111001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4109] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4110] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4111] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4112] = 32'b11000010110001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4113] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4114] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4115] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4116] = 32'b11000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4117] = 32'b01000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4118] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4119] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4120] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4121] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4122] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4123] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4124] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4125] = 32'b11000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4126] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4127] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4128] = 32'b01000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4129] = 32'b11000010111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4130] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4131] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4132] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4133] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4134] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4135] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4136] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4137] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4138] = 32'b11000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4139] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4140] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4141] = 32'b11000011000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4142] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4143] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4144] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4145] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4146] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4147] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4148] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4149] = 32'b11000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4150] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4151] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4152] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4153] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4154] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4155] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4156] = 32'b01000010110001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4157] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4158] = 32'b01000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4159] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4160] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4161] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4162] = 32'b01000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4163] = 32'b11000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4164] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4165] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4166] = 32'b01000010111001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4167] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4168] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4169] = 32'b11000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4170] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4171] = 32'b11000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4172] = 32'b01000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4173] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4174] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4175] = 32'b11000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4176] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4177] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4178] = 32'b01000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4179] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4180] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4181] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4182] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4183] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4184] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4185] = 32'b01000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4186] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4187] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4188] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4189] = 32'b01000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4190] = 32'b11000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4191] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4192] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4193] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4194] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4195] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4196] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4197] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4198] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4199] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4200] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4201] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4202] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4203] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4204] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4205] = 32'b11000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4206] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4207] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4208] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4209] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4210] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4211] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4212] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4213] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4214] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4215] = 32'b01000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4216] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4217] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4218] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4219] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4220] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4221] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4222] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4223] = 32'b01000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4224] = 32'b01000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4225] = 32'b01000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4226] = 32'b01000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4227] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4228] = 32'b01000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4229] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4230] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4231] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4232] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4233] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4234] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4235] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4236] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4237] = 32'b11000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4238] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4239] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4240] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4241] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4242] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4243] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4244] = 32'b11000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4245] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4246] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4247] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4248] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4249] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4250] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4251] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4252] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4253] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4254] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4255] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4256] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4257] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4258] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4259] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4260] = 32'b11000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4261] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4262] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4263] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4264] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4265] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4266] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4267] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4268] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4269] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4270] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4271] = 32'b11000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4272] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4273] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4274] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4275] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4276] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4277] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4278] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4279] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4280] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4281] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4282] = 32'b01000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4283] = 32'b11000010110111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4284] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4285] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4286] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4287] = 32'b01000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4288] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4289] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4290] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4291] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4292] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4293] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4294] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4295] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4296] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4297] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4298] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4299] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4300] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4301] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4302] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4303] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4304] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4305] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4306] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4307] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4308] = 32'b11000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4309] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4310] = 32'b01000010110101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4311] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4312] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4313] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4314] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4315] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4316] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4317] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4318] = 32'b01000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4319] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4320] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4321] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4322] = 32'b01000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4323] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4324] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4325] = 32'b01000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4326] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4327] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4328] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4329] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4330] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4331] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4332] = 32'b11000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4333] = 32'b01000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4334] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4335] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4336] = 32'b01000010110101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4337] = 32'b11000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4338] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4339] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4340] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4341] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4342] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4343] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4344] = 32'b11000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4345] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4346] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4347] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4348] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4349] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4350] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4351] = 32'b11000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4352] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4353] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4354] = 32'b01000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4355] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4356] = 32'b11000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4357] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4358] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4359] = 32'b01000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4360] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4361] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4362] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4363] = 32'b01000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4364] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4365] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4366] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4367] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4368] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4369] = 32'b11000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4370] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4371] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4372] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4373] = 32'b01000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4374] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4375] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4376] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4377] = 32'b01000010110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4378] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4379] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4380] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4381] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4382] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4383] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4384] = 32'b01000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4385] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4386] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4387] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4388] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4389] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4390] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4391] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4392] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4393] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4394] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4395] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4396] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4397] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4398] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4399] = 32'b11000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4400] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4401] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4402] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4403] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4404] = 32'b01000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4405] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4406] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4407] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4408] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4409] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4410] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4411] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4412] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4413] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4414] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4415] = 32'b11000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4416] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4417] = 32'b11000011000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4418] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4419] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4420] = 32'b01000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4421] = 32'b11000010101100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4422] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4423] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4424] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4425] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4426] = 32'b11000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4427] = 32'b11000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4428] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4429] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4430] = 32'b11000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4431] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4432] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4433] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4434] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4435] = 32'b11000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4436] = 32'b01000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4437] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4438] = 32'b11000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4439] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4440] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4441] = 32'b11000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4442] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4443] = 32'b01000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4444] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4445] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4446] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4447] = 32'b11000011000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4448] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4449] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4450] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4451] = 32'b11000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4452] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4453] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4454] = 32'b01000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4455] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4456] = 32'b11000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4457] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4458] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4459] = 32'b11000011000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4460] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4461] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4462] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4463] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4464] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4465] = 32'b11000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4466] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4467] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4468] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4469] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4470] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4471] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4472] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4473] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4474] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4475] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4476] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4477] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4478] = 32'b11000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4479] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4480] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4481] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4482] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4483] = 32'b01000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4484] = 32'b11000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4485] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4486] = 32'b11000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4487] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4488] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4489] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4490] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4491] = 32'b01000010110101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4492] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4493] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4494] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4495] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4496] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4497] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4498] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4499] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4500] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4501] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4502] = 32'b01000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4503] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4504] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4505] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4506] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4507] = 32'b11000010111001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4508] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4509] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4510] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4511] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4512] = 32'b01000010110100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4513] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4514] = 32'b01000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4515] = 32'b01000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4516] = 32'b11000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4517] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4518] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4519] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4520] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4521] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4522] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4523] = 32'b11000010110001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4524] = 32'b01000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4525] = 32'b11000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4526] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4527] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4528] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4529] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4530] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4531] = 32'b01000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4532] = 32'b11000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4533] = 32'b01000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4534] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4535] = 32'b11000010110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4536] = 32'b11000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4537] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4538] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4539] = 32'b01000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4540] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4541] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4542] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4543] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4544] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4545] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4546] = 32'b11000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4547] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4548] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4549] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4550] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4551] = 32'b11000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4552] = 32'b01000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4553] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4554] = 32'b11000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4555] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4556] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4557] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4558] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4559] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4560] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4561] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4562] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4563] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4564] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4565] = 32'b01000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4566] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4567] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4568] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4569] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4570] = 32'b01000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4571] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4572] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4573] = 32'b01000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4574] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4575] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4576] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4577] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4578] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4579] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4580] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4581] = 32'b01000010110111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4582] = 32'b01000010110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4583] = 32'b11000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4584] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4585] = 32'b11000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4586] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4587] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4588] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4589] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4590] = 32'b01000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4591] = 32'b11000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4592] = 32'b01000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4593] = 32'b01000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4594] = 32'b11000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4595] = 32'b11000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4596] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4597] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4598] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4599] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4600] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4601] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4602] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4603] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4604] = 32'b01000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4605] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4606] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4607] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4608] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4609] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4610] = 32'b11000010111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4611] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4612] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4613] = 32'b11000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4614] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4615] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4616] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4617] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4618] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4619] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4620] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4621] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4622] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4623] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4624] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4625] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4626] = 32'b01000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4627] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4628] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4629] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4630] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4631] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4632] = 32'b01000010110011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4633] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4634] = 32'b11000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4635] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4636] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4637] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4638] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4639] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4640] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4641] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4642] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4643] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4644] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4645] = 32'b01000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4646] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4647] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4648] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4649] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4650] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4651] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4652] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4653] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4654] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4655] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4656] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4657] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4658] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4659] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4660] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4661] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4662] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4663] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4664] = 32'b11000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4665] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4666] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4667] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4668] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4669] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4670] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4671] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4672] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4673] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4674] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4675] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4676] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4677] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4678] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4679] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4680] = 32'b11000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4681] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4682] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4683] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4684] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4685] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4686] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4687] = 32'b11000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4688] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4689] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4690] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4691] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4692] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4693] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4694] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4695] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4696] = 32'b11000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4697] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4698] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4699] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4700] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4701] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4702] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4703] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4704] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4705] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4706] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4707] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4708] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4709] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4710] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4711] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4712] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4713] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4714] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4715] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4716] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4717] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4718] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4719] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4720] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4721] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4722] = 32'b11000010110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4723] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4724] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4725] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4726] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4727] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4728] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4729] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4730] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4731] = 32'b11000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4732] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4733] = 32'b01000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4734] = 32'b11000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4735] = 32'b01000010101110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4736] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4737] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4738] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4739] = 32'b11000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4740] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4741] = 32'b11000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4742] = 32'b11000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4743] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4744] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4745] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4746] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4747] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4748] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4749] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4750] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4751] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4752] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4753] = 32'b11000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4754] = 32'b01000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4755] = 32'b01000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4756] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4757] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4758] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4759] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4760] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4761] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4762] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4763] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4764] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4765] = 32'b01000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4766] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4767] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4768] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4769] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4770] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4771] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4772] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4773] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4774] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4775] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4776] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4777] = 32'b11000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4778] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4779] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4780] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4781] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4782] = 32'b01000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4783] = 32'b11000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4784] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4785] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4786] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4787] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4788] = 32'b01000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4789] = 32'b01000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4790] = 32'b01000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4791] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4792] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4793] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4794] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4795] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4796] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4797] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4798] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4799] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4800] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4801] = 32'b01000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4802] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4803] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4804] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4805] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4806] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4807] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4808] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4809] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4810] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4811] = 32'b11000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4812] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4813] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4814] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4815] = 32'b01000010110001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4816] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4817] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4818] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4819] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4820] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4821] = 32'b01000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4822] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4823] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4824] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4825] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4826] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4827] = 32'b11000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4828] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4829] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4830] = 32'b11000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4831] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4832] = 32'b01000010101100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4833] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4834] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4835] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4836] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4837] = 32'b01000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4838] = 32'b11000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4839] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4840] = 32'b11000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4841] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4842] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4843] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4844] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4845] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4846] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4847] = 32'b01000010101100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4848] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4849] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4850] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4851] = 32'b01000010101110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4852] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4853] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4854] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4855] = 32'b01000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4856] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4857] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4858] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4859] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4860] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4861] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4862] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4863] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4864] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4865] = 32'b01000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4866] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4867] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4868] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4869] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4870] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4871] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4872] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4873] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4874] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4875] = 32'b11000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4876] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4877] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4878] = 32'b01000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4879] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4880] = 32'b01000010110001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4881] = 32'b11000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4882] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4883] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4884] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4885] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4886] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4887] = 32'b01000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4888] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4889] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4890] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4891] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4892] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4893] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4894] = 32'b01000010110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4895] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4896] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4897] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4898] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4899] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4900] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4901] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4902] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4903] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4904] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4905] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4906] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4907] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4908] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4909] = 32'b01000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4910] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4911] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4912] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4913] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4914] = 32'b01000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4915] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4916] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4917] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4918] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4919] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4920] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4921] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4922] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4923] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4924] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4925] = 32'b11000010101110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4926] = 32'b01000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4927] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4928] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4929] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4930] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4931] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4932] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4933] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4934] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4935] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4936] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4937] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4938] = 32'b01000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4939] = 32'b11000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4940] = 32'b01000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4941] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4942] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4943] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4944] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4945] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4946] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4947] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4948] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4949] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4950] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4951] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4952] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4953] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4954] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4955] = 32'b01000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4956] = 32'b01000010101100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4957] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4958] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4959] = 32'b11000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4960] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4961] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4962] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4963] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4964] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4965] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4966] = 32'b01000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4967] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4968] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4969] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4970] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4971] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4972] = 32'b11000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4973] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4974] = 32'b01000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4975] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4976] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4977] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4978] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4979] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4980] = 32'b11000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4981] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4982] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4983] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4984] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4985] = 32'b11000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4986] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4987] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4988] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4989] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4990] = 32'b01000010110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4991] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4992] = 32'b11000010101100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4993] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4994] = 32'b11000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4995] = 32'b11000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4996] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4997] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4998] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 4999] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5000] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5001] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5002] = 32'b01000010111001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5003] = 32'b11000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5004] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5005] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5006] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5007] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5008] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5009] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5010] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5011] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5012] = 32'b11000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5013] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5014] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5015] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5016] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5017] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5018] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5019] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5020] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5021] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5022] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5023] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5024] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5025] = 32'b11000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5026] = 32'b11000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5027] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5028] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5029] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5030] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5031] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5032] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5033] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5034] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5035] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5036] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5037] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5038] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5039] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5040] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5041] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5042] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5043] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5044] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5045] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5046] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5047] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5048] = 32'b11000010101110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5049] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5050] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5051] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5052] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5053] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5054] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5055] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5056] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5057] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5058] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5059] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5060] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5061] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5062] = 32'b11000010110001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5063] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5064] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5065] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5066] = 32'b11000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5067] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5068] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5069] = 32'b01000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5070] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5071] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5072] = 32'b11000010110111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5073] = 32'b11000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5074] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5075] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5076] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5077] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5078] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5079] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5080] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5081] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5082] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5083] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5084] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5085] = 32'b01000010101110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5086] = 32'b11000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5087] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5088] = 32'b01000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5089] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5090] = 32'b01000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5091] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5092] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5093] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5094] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5095] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5096] = 32'b11000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5097] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5098] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5099] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5100] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5101] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5102] = 32'b01000010110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5103] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5104] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5105] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5106] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5107] = 32'b01000010110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5108] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5109] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5110] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5111] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5112] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5113] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5114] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5115] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5116] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5117] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5118] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5119] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5120] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5121] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5122] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5123] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5124] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5125] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5126] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5127] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5128] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5129] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5130] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5131] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5132] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5133] = 32'b01000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5134] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5135] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5136] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5137] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5138] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5139] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5140] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5141] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5142] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5143] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5144] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5145] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5146] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5147] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5148] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5149] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5150] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5151] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5152] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5153] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5154] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5155] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5156] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5157] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5158] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5159] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5160] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5161] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5162] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5163] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5164] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5165] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5166] = 32'b11000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5167] = 32'b01000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5168] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5169] = 32'b01000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5170] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5171] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5172] = 32'b11000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5173] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5174] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5175] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5176] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5177] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5178] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5179] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5180] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5181] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5182] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5183] = 32'b11000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5184] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5185] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5186] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5187] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5188] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5189] = 32'b01000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5190] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5191] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5192] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5193] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5194] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5195] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5196] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5197] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5198] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5199] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5200] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5201] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5202] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5203] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5204] = 32'b01000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5205] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5206] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5207] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5208] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5209] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5210] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5211] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5212] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5213] = 32'b11000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5214] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5215] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5216] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5217] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5218] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5219] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5220] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5221] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5222] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5223] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5224] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5225] = 32'b11000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5226] = 32'b01000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5227] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5228] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5229] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5230] = 32'b01000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5231] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5232] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5233] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5234] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5235] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5236] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5237] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5238] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5239] = 32'b11000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5240] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5241] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5242] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5243] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5244] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5245] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5246] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5247] = 32'b01000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5248] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5249] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5250] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5251] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5252] = 32'b11000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5253] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5254] = 32'b11000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5255] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5256] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5257] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5258] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5259] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5260] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5261] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5262] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5263] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5264] = 32'b01000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5265] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5266] = 32'b01000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5267] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5268] = 32'b11000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5269] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5270] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5271] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5272] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5273] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5274] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5275] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5276] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5277] = 32'b01000010110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5278] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5279] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5280] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5281] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5282] = 32'b01000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5283] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5284] = 32'b11000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5285] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5286] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5287] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5288] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5289] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5290] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5291] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5292] = 32'b01000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5293] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5294] = 32'b11000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5295] = 32'b11000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5296] = 32'b01000010110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5297] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5298] = 32'b01000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5299] = 32'b11000010110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5300] = 32'b11000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5301] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5302] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5303] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5304] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5305] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5306] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5307] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5308] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5309] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5310] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5311] = 32'b11000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5312] = 32'b01000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5313] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5314] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5315] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5316] = 32'b01000010110001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5317] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5318] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5319] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5320] = 32'b11000010110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5321] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5322] = 32'b11000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5323] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5324] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5325] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5326] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5327] = 32'b01000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5328] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5329] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5330] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5331] = 32'b01000010111001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5332] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5333] = 32'b01000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5334] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5335] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5336] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5337] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5338] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5339] = 32'b11000010110100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5340] = 32'b01000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5341] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5342] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5343] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5344] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5345] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5346] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5347] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5348] = 32'b11000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5349] = 32'b01000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5350] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5351] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5352] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5353] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5354] = 32'b01000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5355] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5356] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5357] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5358] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5359] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5360] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5361] = 32'b01000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5362] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5363] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5364] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5365] = 32'b11000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5366] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5367] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5368] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5369] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5370] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5371] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5372] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5373] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5374] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5375] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5376] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5377] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5378] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5379] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5380] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5381] = 32'b01000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5382] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5383] = 32'b11000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5384] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5385] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5386] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5387] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5388] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5389] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5390] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5391] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5392] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5393] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5394] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5395] = 32'b11000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5396] = 32'b01000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5397] = 32'b01000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5398] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5399] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5400] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5401] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5402] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5403] = 32'b01000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5404] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5405] = 32'b01000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5406] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5407] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5408] = 32'b11000010101110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5409] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5410] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5411] = 32'b11000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5412] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5413] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5414] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5415] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5416] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5417] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5418] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5419] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5420] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5421] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5422] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5423] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5424] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5425] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5426] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5427] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5428] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5429] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5430] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5431] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5432] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5433] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5434] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5435] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5436] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5437] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5438] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5439] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5440] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5441] = 32'b11000010110101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5442] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5443] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5444] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5445] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5446] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5447] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5448] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5449] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5450] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5451] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5452] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5453] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5454] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5455] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5456] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5457] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5458] = 32'b11000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5459] = 32'b11000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5460] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5461] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5462] = 32'b11000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5463] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5464] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5465] = 32'b11000011000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5466] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5467] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5468] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5469] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5470] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5471] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5472] = 32'b01000010111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5473] = 32'b01000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5474] = 32'b01000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5475] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5476] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5477] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5478] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5479] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5480] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5481] = 32'b01000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5482] = 32'b11000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5483] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5484] = 32'b01000010101110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5485] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5486] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5487] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5488] = 32'b01000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5489] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5490] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5491] = 32'b11000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5492] = 32'b01000010110100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5493] = 32'b11000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5494] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5495] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5496] = 32'b01000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5497] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5498] = 32'b11000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5499] = 32'b01000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5500] = 32'b01000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5501] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5502] = 32'b01000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5503] = 32'b01000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5504] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5505] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5506] = 32'b11000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5507] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5508] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5509] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5510] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5511] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5512] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5513] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5514] = 32'b01000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5515] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5516] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5517] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5518] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5519] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5520] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5521] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5522] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5523] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5524] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5525] = 32'b11000010101110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5526] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5527] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5528] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5529] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5530] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5531] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5532] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5533] = 32'b11000011000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5534] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5535] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5536] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5537] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5538] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5539] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5540] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5541] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5542] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5543] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5544] = 32'b01000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5545] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5546] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5547] = 32'b11000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5548] = 32'b11000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5549] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5550] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5551] = 32'b01000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5552] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5553] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5554] = 32'b11000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5555] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5556] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5557] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5558] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5559] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5560] = 32'b11000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5561] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5562] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5563] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5564] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5565] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5566] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5567] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5568] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5569] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5570] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5571] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5572] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5573] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5574] = 32'b11000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5575] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5576] = 32'b01000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5577] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5578] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5579] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5580] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5581] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5582] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5583] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5584] = 32'b11000010110100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5585] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5586] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5587] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5588] = 32'b11000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5589] = 32'b01000010101100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5590] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5591] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5592] = 32'b11000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5593] = 32'b01000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5594] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5595] = 32'b01000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5596] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5597] = 32'b01000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5598] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5599] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5600] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5601] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5602] = 32'b11000011000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5603] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5604] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5605] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5606] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5607] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5608] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5609] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5610] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5611] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5612] = 32'b11000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5613] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5614] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5615] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5616] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5617] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5618] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5619] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5620] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5621] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5622] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5623] = 32'b11000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5624] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5625] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5626] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5627] = 32'b01000010101110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5628] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5629] = 32'b01000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5630] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5631] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5632] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5633] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5634] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5635] = 32'b11000011000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5636] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5637] = 32'b01000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5638] = 32'b11000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5639] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5640] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5641] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5642] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5643] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5644] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5645] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5646] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5647] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5648] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5649] = 32'b11000010110111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5650] = 32'b01000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5651] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5652] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5653] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5654] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5655] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5656] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5657] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5658] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5659] = 32'b11000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5660] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5661] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5662] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5663] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5664] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5665] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5666] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5667] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5668] = 32'b01000010110101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5669] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5670] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5671] = 32'b11000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5672] = 32'b01000010110100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5673] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5674] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5675] = 32'b01000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5676] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5677] = 32'b11000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5678] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5679] = 32'b01000010110001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5680] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5681] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5682] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5683] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5684] = 32'b01000010101100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5685] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5686] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5687] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5688] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5689] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5690] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5691] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5692] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5693] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5694] = 32'b11000010110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5695] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5696] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5697] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5698] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5699] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5700] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5701] = 32'b11000010110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5702] = 32'b01000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5703] = 32'b11000010111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5704] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5705] = 32'b11000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5706] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5707] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5708] = 32'b01000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5709] = 32'b11000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5710] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5711] = 32'b01000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5712] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5713] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5714] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5715] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5716] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5717] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5718] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5719] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5720] = 32'b11000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5721] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5722] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5723] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5724] = 32'b11000010110001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5725] = 32'b11000010110111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5726] = 32'b01000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5727] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5728] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5729] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5730] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5731] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5732] = 32'b11000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5733] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5734] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5735] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5736] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5737] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5738] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5739] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5740] = 32'b01000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5741] = 32'b11000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5742] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5743] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5744] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5745] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5746] = 32'b11000010110101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5747] = 32'b11000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5748] = 32'b11000010111011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5749] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5750] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5751] = 32'b11000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5752] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5753] = 32'b01000010110100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5754] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5755] = 32'b01000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5756] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5757] = 32'b01000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5758] = 32'b01000010111001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5759] = 32'b11000011000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5760] = 32'b11000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5761] = 32'b11000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5762] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5763] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5764] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5765] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5766] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5767] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5768] = 32'b11000010100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5769] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5770] = 32'b11000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5771] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5772] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5773] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5774] = 32'b11000010100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5775] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5776] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5777] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5778] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5779] = 32'b11000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5780] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5781] = 32'b11000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5782] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5783] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5784] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5785] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5786] = 32'b11000010110101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5787] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5788] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5789] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5790] = 32'b11000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5791] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5792] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5793] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5794] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5795] = 32'b11000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5796] = 32'b11000010110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5797] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5798] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5799] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5800] = 32'b11000010110011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5801] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5802] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5803] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5804] = 32'b11000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5805] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5806] = 32'b11000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5807] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5808] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5809] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5810] = 32'b01000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5811] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5812] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5813] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5814] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5815] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5816] = 32'b01000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5817] = 32'b01000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5818] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5819] = 32'b01000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5820] = 32'b01000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5821] = 32'b01000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5822] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5823] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5824] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5825] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5826] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5827] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5828] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5829] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5830] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5831] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5832] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5833] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5834] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5835] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5836] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5837] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5838] = 32'b01000010110011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5839] = 32'b01000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5840] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5841] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5842] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5843] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5844] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5845] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5846] = 32'b11000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5847] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5848] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5849] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5850] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5851] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5852] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5853] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5854] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5855] = 32'b01000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5856] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5857] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5858] = 32'b11000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5859] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5860] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5861] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5862] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5863] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5864] = 32'b01000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5865] = 32'b01000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5866] = 32'b11000010110101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5867] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5868] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5869] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5870] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5871] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5872] = 32'b01000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5873] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5874] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5875] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5876] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5877] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5878] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5879] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5880] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5881] = 32'b11000010110011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5882] = 32'b01000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5883] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5884] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5885] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5886] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5887] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5888] = 32'b01000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5889] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5890] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5891] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5892] = 32'b01000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5893] = 32'b01000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5894] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5895] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5896] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5897] = 32'b01000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5898] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5899] = 32'b01000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5900] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5901] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5902] = 32'b01000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5903] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5904] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5905] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5906] = 32'b01000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5907] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5908] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5909] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5910] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5911] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5912] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5913] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5914] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5915] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5916] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5917] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5918] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5919] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5920] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5921] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5922] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5923] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5924] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5925] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5926] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5927] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5928] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5929] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5930] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5931] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5932] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5933] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5934] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5935] = 32'b11000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5936] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5937] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5938] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5939] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5940] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5941] = 32'b01000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5942] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5943] = 32'b11000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5944] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5945] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5946] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5947] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5948] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5949] = 32'b01000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5950] = 32'b11000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5951] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5952] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5953] = 32'b01000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5954] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5955] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5956] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5957] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5958] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5959] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5960] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5961] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5962] = 32'b11000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5963] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5964] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5965] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5966] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5967] = 32'b11000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5968] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5969] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5970] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5971] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5972] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5973] = 32'b11000010101110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5974] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5975] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5976] = 32'b11000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5977] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5978] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5979] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5980] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5981] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5982] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5983] = 32'b01000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5984] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5985] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5986] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5987] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5988] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5989] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5990] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5991] = 32'b11000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5992] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5993] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5994] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5995] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5996] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5997] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5998] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 5999] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6000] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6001] = 32'b11000010110100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6002] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6003] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6004] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6005] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6006] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6007] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6008] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6009] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6010] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6011] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6012] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6013] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6014] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6015] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6016] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6017] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6018] = 32'b11000010110100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6019] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6020] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6021] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6022] = 32'b11000010111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6023] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6024] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6025] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6026] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6027] = 32'b01000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6028] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6029] = 32'b01000010110100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6030] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6031] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6032] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6033] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6034] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6035] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6036] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6037] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6038] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6039] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6040] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6041] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6042] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6043] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6044] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6045] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6046] = 32'b11000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6047] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6048] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6049] = 32'b01000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6050] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6051] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6052] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6053] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6054] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6055] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6056] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6057] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6058] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6059] = 32'b11000010110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6060] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6061] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6062] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6063] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6064] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6065] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6066] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6067] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6068] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6069] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6070] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6071] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6072] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6073] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6074] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6075] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6076] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6077] = 32'b01000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6078] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6079] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6080] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6081] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6082] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6083] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6084] = 32'b11000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6085] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6086] = 32'b01000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6087] = 32'b01000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6088] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6089] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6090] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6091] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6092] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6093] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6094] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6095] = 32'b01000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6096] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6097] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6098] = 32'b01000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6099] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6100] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6101] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6102] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6103] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6104] = 32'b11000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6105] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6106] = 32'b11000010110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6107] = 32'b01000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6108] = 32'b01000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6109] = 32'b01000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6110] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6111] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6112] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6113] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6114] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6115] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6116] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6117] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6118] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6119] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6120] = 32'b01000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6121] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6122] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6123] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6124] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6125] = 32'b01000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6126] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6127] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6128] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6129] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6130] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6131] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6132] = 32'b01000010110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6133] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6134] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6135] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6136] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6137] = 32'b01000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6138] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6139] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6140] = 32'b11000010110001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6141] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6142] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6143] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6144] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6145] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6146] = 32'b11000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6147] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6148] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6149] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6150] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6151] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6152] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6153] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6154] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6155] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6156] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6157] = 32'b11000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6158] = 32'b01000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6159] = 32'b11000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6160] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6161] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6162] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6163] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6164] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6165] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6166] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6167] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6168] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6169] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6170] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6171] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6172] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6173] = 32'b01000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6174] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6175] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6176] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6177] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6178] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6179] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6180] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6181] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6182] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6183] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6184] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6185] = 32'b11000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6186] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6187] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6188] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6189] = 32'b11000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6190] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6191] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6192] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6193] = 32'b11000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6194] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6195] = 32'b01000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6196] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6197] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6198] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6199] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6200] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6201] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6202] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6203] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6204] = 32'b11000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6205] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6206] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6207] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6208] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6209] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6210] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6211] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6212] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6213] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6214] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6215] = 32'b01000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6216] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6217] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6218] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6219] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6220] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6221] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6222] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6223] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6224] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6225] = 32'b11000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6226] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6227] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6228] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6229] = 32'b11000010110101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6230] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6231] = 32'b01000010110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6232] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6233] = 32'b01000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6234] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6235] = 32'b11000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6236] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6237] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6238] = 32'b11000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6239] = 32'b01000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6240] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6241] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6242] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6243] = 32'b11000010101110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6244] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6245] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6246] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6247] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6248] = 32'b11000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6249] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6250] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6251] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6252] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6253] = 32'b01000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6254] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6255] = 32'b01000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6256] = 32'b01000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6257] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6258] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6259] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6260] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6261] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6262] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6263] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6264] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6265] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6266] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6267] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6268] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6269] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6270] = 32'b01000010111001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6271] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6272] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6273] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6274] = 32'b11000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6275] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6276] = 32'b11000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6277] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6278] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6279] = 32'b01000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6280] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6281] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6282] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6283] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6284] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6285] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6286] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6287] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6288] = 32'b11000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6289] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6290] = 32'b11000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6291] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6292] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6293] = 32'b01000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6294] = 32'b11000010110111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6295] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6296] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6297] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6298] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6299] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6300] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6301] = 32'b11000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6302] = 32'b11000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6303] = 32'b11000010110101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6304] = 32'b01000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6305] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6306] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6307] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6308] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6309] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6310] = 32'b11000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6311] = 32'b01000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6312] = 32'b01000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6313] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6314] = 32'b11000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6315] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6316] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6317] = 32'b01000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6318] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6319] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6320] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6321] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6322] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6323] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6324] = 32'b11000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6325] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6326] = 32'b01000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6327] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6328] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6329] = 32'b01000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6330] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6331] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6332] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6333] = 32'b01000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6334] = 32'b11000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6335] = 32'b11000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6336] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6337] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6338] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6339] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6340] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6341] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6342] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6343] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6344] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6345] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6346] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6347] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6348] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6349] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6350] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6351] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6352] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6353] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6354] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6355] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6356] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6357] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6358] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6359] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6360] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6361] = 32'b11000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6362] = 32'b11000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6363] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6364] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6365] = 32'b11000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6366] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6367] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6368] = 32'b01000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6369] = 32'b11000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6370] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6371] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6372] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6373] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6374] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6375] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6376] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6377] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6378] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6379] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6380] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6381] = 32'b11000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6382] = 32'b11000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6383] = 32'b11000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6384] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6385] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6386] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6387] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6388] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6389] = 32'b11000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6390] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6391] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6392] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6393] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6394] = 32'b11000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6395] = 32'b01000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6396] = 32'b11000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6397] = 32'b01000010110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6398] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6399] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6400] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6401] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6402] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6403] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6404] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6405] = 32'b01000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6406] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6407] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6408] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6409] = 32'b11000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6410] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6411] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6412] = 32'b01000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6413] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6414] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6415] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6416] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6417] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6418] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6419] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6420] = 32'b11000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6421] = 32'b11000010010111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6422] = 32'b01000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6423] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6424] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6425] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6426] = 32'b11000010110111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6427] = 32'b01000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6428] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6429] = 32'b11000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6430] = 32'b01000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6431] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6432] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6433] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6434] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6435] = 32'b01000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6436] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6437] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6438] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6439] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6440] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6441] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6442] = 32'b01000010111001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6443] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6444] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6445] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6446] = 32'b01000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6447] = 32'b11000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6448] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6449] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6450] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6451] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6452] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6453] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6454] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6455] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6456] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6457] = 32'b01000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6458] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6459] = 32'b11000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6460] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6461] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6462] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6463] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6464] = 32'b01000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6465] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6466] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6467] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6468] = 32'b11000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6469] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6470] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6471] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6472] = 32'b01000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6473] = 32'b11000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6474] = 32'b01000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6475] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6476] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6477] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6478] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6479] = 32'b01000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6480] = 32'b11000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6481] = 32'b11000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6482] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6483] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6484] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6485] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6486] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6487] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6488] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6489] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6490] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6491] = 32'b01000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6492] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6493] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6494] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6495] = 32'b01000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6496] = 32'b01000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6497] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6498] = 32'b01000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6499] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6500] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6501] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6502] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6503] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6504] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6505] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6506] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6507] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6508] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6509] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6510] = 32'b01000010101100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6511] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6512] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6513] = 32'b01000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6514] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6515] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6516] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6517] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6518] = 32'b01000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6519] = 32'b01000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6520] = 32'b01000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6521] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6522] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6523] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6524] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6525] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6526] = 32'b01000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6527] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6528] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6529] = 32'b01000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6530] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6531] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6532] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6533] = 32'b01000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6534] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6535] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6536] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6537] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6538] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6539] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6540] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6541] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6542] = 32'b01000010110011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6543] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6544] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6545] = 32'b01000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6546] = 32'b11000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6547] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6548] = 32'b01000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6549] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6550] = 32'b11000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6551] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6552] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6553] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6554] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6555] = 32'b11000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6556] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6557] = 32'b01000010110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6558] = 32'b11000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6559] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6560] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6561] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6562] = 32'b01000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6563] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6564] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6565] = 32'b01000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6566] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6567] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6568] = 32'b11000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6569] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6570] = 32'b01000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6571] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6572] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6573] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6574] = 32'b11000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6575] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6576] = 32'b01000010111110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6577] = 32'b11000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6578] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6579] = 32'b01000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6580] = 32'b11000010001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6581] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6582] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6583] = 32'b11000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6584] = 32'b01000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6585] = 32'b11000010010010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6586] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6587] = 32'b11000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6588] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6589] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6590] = 32'b11000010101111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6591] = 32'b01000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6592] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6593] = 32'b11000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6594] = 32'b11000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6595] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6596] = 32'b11000010010110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6597] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6598] = 32'b01000010100011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6599] = 32'b11000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6600] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6601] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6602] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6603] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6604] = 32'b11000010110001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6605] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6606] = 32'b01000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6607] = 32'b11000010110110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6608] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6609] = 32'b11000010100010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6610] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6611] = 32'b11000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6612] = 32'b11000010110111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6613] = 32'b11000010011011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6614] = 32'b00111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6615] = 32'b01000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6616] = 32'b11000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6617] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6618] = 32'b01000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6619] = 32'b01000010110011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6620] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6621] = 32'b11000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6622] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6623] = 32'b01000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6624] = 32'b01000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6625] = 32'b11000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6626] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6627] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6628] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6629] = 32'b01000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6630] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6631] = 32'b11000010110101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6632] = 32'b11000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6633] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6634] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6635] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6636] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6637] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6638] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6639] = 32'b01000010000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6640] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6641] = 32'b01000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6642] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6643] = 32'b11000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6644] = 32'b11000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6645] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6646] = 32'b11000010101001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6647] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6648] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6649] = 32'b11000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6650] = 32'b11000010101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6651] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6652] = 32'b01000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6653] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6654] = 32'b01000000110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6655] = 32'b01000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6656] = 32'b11000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6657] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6658] = 32'b01000010011010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6659] = 32'b11000010100110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6660] = 32'b11000001110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6661] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6662] = 32'b01000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6663] = 32'b01000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6664] = 32'b01000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6665] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6666] = 32'b01000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6667] = 32'b11000010111000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6668] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6669] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6670] = 32'b11000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6671] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6672] = 32'b11000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6673] = 32'b11000010111001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6674] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6675] = 32'b11000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6676] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6677] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6678] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6679] = 32'b11000010111101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6680] = 32'b01000010110111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6681] = 32'b01000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6682] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6683] = 32'b11000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6684] = 32'b01000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6685] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6686] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6687] = 32'b01000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6688] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6689] = 32'b11000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6690] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6691] = 32'b11000010101101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6692] = 32'b11000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6693] = 32'b01000010010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6694] = 32'b01000010100000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6695] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6696] = 32'b11000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6697] = 32'b01000010101110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6698] = 32'b01000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6699] = 32'b11000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6700] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6701] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6702] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6703] = 32'b11000010100111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6704] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6705] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6706] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6707] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6708] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6709] = 32'b01000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6710] = 32'b11000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6711] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6712] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6713] = 32'b01000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6714] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6715] = 32'b01000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6716] = 32'b11000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6717] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6718] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6719] = 32'b11000010111101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6720] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6721] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6722] = 32'b11000010101111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6723] = 32'b01000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6724] = 32'b01000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6725] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6726] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6727] = 32'b11000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6728] = 32'b01000010011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6729] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6730] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6731] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6732] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6733] = 32'b11000001100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6734] = 32'b11000010111010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6735] = 32'b11000010110101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6736] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6737] = 32'b11000010110001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6738] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6739] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6740] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6741] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6742] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6743] = 32'b11000010110010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6744] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6745] = 32'b11000010101001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6746] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6747] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6748] = 32'b01000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6749] = 32'b01000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6750] = 32'b01000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6751] = 32'b01000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6752] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6753] = 32'b11000010011001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6754] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6755] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6756] = 32'b01000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6757] = 32'b11000001000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6758] = 32'b11000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6759] = 32'b11000010100101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6760] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6761] = 32'b11000010110100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6762] = 32'b01000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6763] = 32'b01000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6764] = 32'b11000010010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6765] = 32'b01000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6766] = 32'b11000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6767] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6768] = 32'b01000000101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6769] = 32'b11000010111111100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6770] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6771] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6772] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6773] = 32'b11000001011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6774] = 32'b01000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6775] = 32'b01000010101110100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6776] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6777] = 32'b00000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6778] = 32'b11000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6779] = 32'b01000010100001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6780] = 32'b01000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6781] = 32'b01000000111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6782] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6783] = 32'b01000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6784] = 32'b01000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6785] = 32'b01000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6786] = 32'b01000010101000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6787] = 32'b01000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6788] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6789] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6790] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6791] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6792] = 32'b01000010010011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6793] = 32'b11000010000111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6794] = 32'b01000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6795] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6796] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6797] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6798] = 32'b01000010011110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6799] = 32'b01000010101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6800] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6801] = 32'b01000010100100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6802] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6803] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6804] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6805] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6806] = 32'b01000010110011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6807] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6808] = 32'b11000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6809] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6810] = 32'b11000010101010100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6811] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6812] = 32'b11000001010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6813] = 32'b01000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6814] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6815] = 32'b11000010101100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6816] = 32'b01000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6817] = 32'b11000001110010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6818] = 32'b01000010111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6819] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6820] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6821] = 32'b01000010011111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6822] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6823] = 32'b01000010011000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6824] = 32'b11000010100001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6825] = 32'b11000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6826] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6827] = 32'b01000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6828] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6829] = 32'b01000010101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6830] = 32'b01000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6831] = 32'b11000010100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6832] = 32'b01000001101110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6833] = 32'b01000001100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6834] = 32'b11000010001110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6835] = 32'b01000010111111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6836] = 32'b01000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6837] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6838] = 32'b11000010010101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6839] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6840] = 32'b01000010101101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6841] = 32'b01000001101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6842] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6843] = 32'b11000010001111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6844] = 32'b11000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6845] = 32'b01000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6846] = 32'b01000001111000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6847] = 32'b11000010100010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6848] = 32'b01000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6849] = 32'b01000010110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6850] = 32'b11000001110000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6851] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6852] = 32'b11000010110000100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6853] = 32'b11000001010100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6854] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6855] = 32'b11000001110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6856] = 32'b11000001101010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6857] = 32'b11000010110100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6858] = 32'b11000001101100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6859] = 32'b11000010011101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6860] = 32'b11000010111011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6861] = 32'b11000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6862] = 32'b11000010001001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6863] = 32'b11000000010000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6864] = 32'b11000010101011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6865] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6866] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6867] = 32'b01000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6868] = 32'b10111111100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6869] = 32'b11000010001010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6870] = 32'b11000000000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6871] = 32'b01000010001101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6872] = 32'b01000010001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6873] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6874] = 32'b11000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6875] = 32'b11000010000110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6876] = 32'b11000010000001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6877] = 32'b11000010000100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6878] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6879] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6880] = 32'b01000010100101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6881] = 32'b01000010110001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6882] = 32'b11000001000000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6883] = 32'b01000010110101100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6884] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6885] = 32'b01000001001100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6886] = 32'b01000010111100100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6887] = 32'b11000001111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6888] = 32'b11000010010001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6889] = 32'b11000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6890] = 32'b11000010000101000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6891] = 32'b01000010001011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6892] = 32'b11000010101000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6893] = 32'b11000001111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6894] = 32'b01000001100110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6895] = 32'b01000001011100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6896] = 32'b01000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6897] = 32'b11000010100011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6898] = 32'b01000010100111000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6899] = 32'b11000010110110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6900] = 32'b11000010101011100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6901] = 32'b01000010000010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6902] = 32'b11000000100000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6903] = 32'b11000001111100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6904] = 32'b11000010110001000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6905] = 32'b01000010111110000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6906] = 32'b11000010111001100000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6907] = 32'b11000001100100000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6908] = 32'b11000010111010000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6909] = 32'b01000010000011000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6910] = 32'b01000001001000000000000000000000;
	assign	noise_gru_recurrent_weights_array[ 6911] = 32'b11000010111110100000000000000000;

}
//////////////////////////////////////////////////////////////////////////////////////////////////
	generate 
		genvar i, bit;
		for ( i = 0 ; i < 144 ; i = i + 1 ) 
			for ( bit = 0 ; bit < 32 ; bit = bit + 1 ) begin	
				assign noise_gru_bias[i*bit] = noise_gru_bias_array[i][bit];	
			end

		for ( i = 0 ; i < 12960 ; i = i + 1 ) 
			for ( bit = 0 ; bit < 32 ; bit = bit + 1 ) begin	
				assign noise_gru_input_weights[i*bit] = noise_gru_input_weights_array[i][bit];	
			end

		for ( i = 0 ; i < 6912 ; i = i + 1 ) 
			for ( bit = 0 ; bit < 32 ; bit = bit + 1 ) begin	
				assign noise_gru_recurrent_weights[i*bit] = noise_gru_recurrent_weights_array[i][bit];	
			end
	endgenerate	


	initial	begin 
		weights_scale	= 32'b0_01110111_00000000000000000000000;  // 1.f/256
		tmpsum1		= 0;
		tmpsum2		= 0;
		z 		= 0;
		r 		= 0;
		h 		= 0;
	end

	always @(posedge clk) begin

		if(index1 < N) begin

			sum	<= noise_gru_bias[index1*float +: float];

			if(index2 < M) begin
				tmpsum1	<= noise_gru_input_weights[(index2*stride+index1)*float +: float] * noise_input[index2*float +: float];
				sum	<= tmpsum1 + sum;
				index2	<= index2 + 1;
			end

			if(index3 < M) begin
				tmpsum2	<= noise_gru_recurrent_weights[(index3*stride+index1)*float +: float] * noise_gru_state[index3*float +: float];
				sum	<= tmpsum2 + sum;
				index3	<= index3 + 1;
			end

			index1	<= index1 + 1;

			tmpz[index1*float +: 32] <= weights_scale * sum;
		end
	end

	sigmoid sigforz(tmpz, z);

	always @(posedge clk) begin

		index1 =0; index2 =0; index3 = 0;

		if(index1 < N) begin

			sum	<= noise_gru_bias[index1*float+N +: 32];

			if(index2 < M) begin
				tmpsum1	<= noise_gru_input_weights[(N+index2*stride+index1)*float +: float] * noise_input[index2*float +: float];
				sum	<= tmpsum1 + sum;
				index2	<= index2 + 1;
			end

			if(index3 < M) begin
				tmpsum2	<= noise_gru_recurrent_weights[(N+index3*stride+index1)*float +: float] * noise_gru_state[index3*float +: float];
				sum	<= tmpsum2 + sum;
				index3	<= index3 + 1;
			end

			index1	<= index1 + 1;

			tmpr[index1*float +: 32] <= weights_scale * sum;
		end
	end
	sigmoid sigforh(tmpr, r);

	always @(posedge clk) begin

		index1 =0; index2 =0; index3 = 0;

		tmpsum1 = 0; tmpsum2 = 0;

		if(index1 < N) begin

			sum	<= noise_gru_bias[2*N+index1*float+N +: 32];

			if(index2 < M) begin
				tmpsum1	<= noise_gru_input_weights[(2*N+index2*stride+index1)*float +: float] * noise_input[index2*float +: float];
				sum	<= tmpsum1 + sum;
				index2	<= index2 + 1;
			end

			if(index3 < M) begin
				tmpsum2	<= noise_gru_recurrent_weights[(2*N+index3*stride+index1)*float +:float] * noise_gru_state[index3*float +: float] * r[index3*float +: float];
				sum	<= tmpsum2 + sum;
				index3	<= index3 + 1;
			end

			// relu reluforg2(sum, tmptmp);

			h[index1*float +: float] = z[index1*float +: float] * noise_gru_state[index1*float +: float] + (one - z[index1*float +: float]) * tmptmp;

			index1	<= index1 + 1;
		end
	end
	
	assign noise_gru_state = h;

endmodule
	