module gru1 ( vad_gru_state, dense_out, clk );	// 24 -> 24

	parameter 			float = 32;

	reg	[          float : 0]	vad_gru_bias_array[71:0];
	wire	[(   72*float)-1 : 0]	vad_gru_bias;

	reg	[          float : 0]	vad_gru_input_weights_array[1727:0];
	wire	[( 1728*float)-1 : 0]	vad_gru_input_weights;

	reg	[          float : 0]	vad_gru_recurrent_weights_array[1727:0];
	wire	[( 1728*float)-1 : 0]	vad_gru_recurrent_weights;


	output 	[(   24*float)-1 : 0]	vad_gru_state;
	input 	[(   24*float)-1 : 0]	dense_out;
	input 							clk;
	
	reg	[(   24*float)-1 : 0]	z ,tmpz, r, tmpr, h, tmph, tmptmp;
	reg	[        float-1 : 0]	weights_scale;
	reg	[(   24*float)-1 : 0]	sum, tmpsum1, tmpsum2;

	integer	index1		= 0;
	integer	index2		= 0;
	integer	index3		= 0;
	integer	M		= 24;
	integer	N		= 24;
	integer	stride		= 72;
	integer	one		= 1;
////////////////////////////////////////////////////////////////////////////////
{
	assign	vad_gru_bias_array[    0] = 32'b01000010111110000000000000000000;
	assign	vad_gru_bias_array[    1] = 32'b01000010111110100000000000000000;
	assign	vad_gru_bias_array[    2] = 32'b11000010011001000000000000000000;
	assign	vad_gru_bias_array[    3] = 32'b11000010111111000000000000000000;
	assign	vad_gru_bias_array[    4] = 32'b01000010010101000000000000000000;
	assign	vad_gru_bias_array[    5] = 32'b01000010111101100000000000000000;
	assign	vad_gru_bias_array[    6] = 32'b01000010111111100000000000000000;
	assign	vad_gru_bias_array[    7] = 32'b11000010100101100000000000000000;
	assign	vad_gru_bias_array[    8] = 32'b01000010100010000000000000000000;
	assign	vad_gru_bias_array[    9] = 32'b01000010110011000000000000000000;
	assign	vad_gru_bias_array[   10] = 32'b11000000000000000000000000000000;
	assign	vad_gru_bias_array[   11] = 32'b01000010111010000000000000000000;
	assign	vad_gru_bias_array[   12] = 32'b01000010111110000000000000000000;
	assign	vad_gru_bias_array[   13] = 32'b01000010111111100000000000000000;
	assign	vad_gru_bias_array[   14] = 32'b01000010111110000000000000000000;
	assign	vad_gru_bias_array[   15] = 32'b01000010111110100000000000000000;
	assign	vad_gru_bias_array[   16] = 32'b01000010111111000000000000000000;
	assign	vad_gru_bias_array[   17] = 32'b01000010111101100000000000000000;
	assign	vad_gru_bias_array[   18] = 32'b11000001100000000000000000000000;
	assign	vad_gru_bias_array[   19] = 32'b01000010010000000000000000000000;
	assign	vad_gru_bias_array[   20] = 32'b01000010111110100000000000000000;
	assign	vad_gru_bias_array[   21] = 32'b01000010111111000000000000000000;
	assign	vad_gru_bias_array[   22] = 32'b01000010100111000000000000000000;
	assign	vad_gru_bias_array[   23] = 32'b01000010101010100000000000000000;
	assign	vad_gru_bias_array[   24] = 32'b01000001001100000000000000000000;
	assign	vad_gru_bias_array[   25] = 32'b01000010111111000000000000000000;
	assign	vad_gru_bias_array[   26] = 32'b11000001111100000000000000000000;
	assign	vad_gru_bias_array[   27] = 32'b11000001111100000000000000000000;
	assign	vad_gru_bias_array[   28] = 32'b11000010100000000000000000000000;
	assign	vad_gru_bias_array[   29] = 32'b11000000010000000000000000000000;
	assign	vad_gru_bias_array[   30] = 32'b11000010110100100000000000000000;
	assign	vad_gru_bias_array[   31] = 32'b11000001111010000000000000000000;
	assign	vad_gru_bias_array[   32] = 32'b11000001100010000000000000000000;
	assign	vad_gru_bias_array[   33] = 32'b01000010100010100000000000000000;
	assign	vad_gru_bias_array[   34] = 32'b01000010011111000000000000000000;
	assign	vad_gru_bias_array[   35] = 32'b01000000000000000000000000000000;
	assign	vad_gru_bias_array[   36] = 32'b11000010000000000000000000000000;
	assign	vad_gru_bias_array[   37] = 32'b11000001001000000000000000000000;
	assign	vad_gru_bias_array[   38] = 32'b11000010011110000000000000000000;
	assign	vad_gru_bias_array[   39] = 32'b01000010111000100000000000000000;
	assign	vad_gru_bias_array[   40] = 32'b11000010010100000000000000000000;
	assign	vad_gru_bias_array[   41] = 32'b01000010111000000000000000000000;
	assign	vad_gru_bias_array[   42] = 32'b11000010110110100000000000000000;
	assign	vad_gru_bias_array[   43] = 32'b01000010111000000000000000000000;
	assign	vad_gru_bias_array[   44] = 32'b01000000111000000000000000000000;
	assign	vad_gru_bias_array[   45] = 32'b11000010001000000000000000000000;
	assign	vad_gru_bias_array[   46] = 32'b01000010100100100000000000000000;
	assign	vad_gru_bias_array[   47] = 32'b01000010010101000000000000000000;
	assign	vad_gru_bias_array[   48] = 32'b01000010011110000000000000000000;
	assign	vad_gru_bias_array[   49] = 32'b01000000110000000000000000000000;
	assign	vad_gru_bias_array[   50] = 32'b11000000000000000000000000000000;
	assign	vad_gru_bias_array[   51] = 32'b00000000000000000000000000000000;
	assign	vad_gru_bias_array[   52] = 32'b00000000000000000000000000000000;
	assign	vad_gru_bias_array[   53] = 32'b01000010110010000000000000000000;
	assign	vad_gru_bias_array[   54] = 32'b11000001100000000000000000000000;
	assign	vad_gru_bias_array[   55] = 32'b01000001110100000000000000000000;
	assign	vad_gru_bias_array[   56] = 32'b11000001110000000000000000000000;
	assign	vad_gru_bias_array[   57] = 32'b01000010011000000000000000000000;
	assign	vad_gru_bias_array[   58] = 32'b01000001110100000000000000000000;
	assign	vad_gru_bias_array[   59] = 32'b11000001001000000000000000000000;
	assign	vad_gru_bias_array[   60] = 32'b11000010000001000000000000000000;
	assign	vad_gru_bias_array[   61] = 32'b01000010001001000000000000000000;
	assign	vad_gru_bias_array[   62] = 32'b01000010100011000000000000000000;
	assign	vad_gru_bias_array[   63] = 32'b01000010110110100000000000000000;
	assign	vad_gru_bias_array[   64] = 32'b11000001111010000000000000000000;
	assign	vad_gru_bias_array[   65] = 32'b01000010111111100000000000000000;
	assign	vad_gru_bias_array[   66] = 32'b01000010000010000000000000000000;
	assign	vad_gru_bias_array[   67] = 32'b11000010100001000000000000000000;
	assign	vad_gru_bias_array[   68] = 32'b01000010010001000000000000000000;
	assign	vad_gru_bias_array[   69] = 32'b01000010010101000000000000000000;
	assign	vad_gru_bias_array[   70] = 32'b01000001110110000000000000000000;
	assign	vad_gru_bias_array[   71] = 32'b01000010011110000000000000000000;

	assign	vad_gru_input_weights_array[    0] = 32'b11000010111110000000000000000000;
	assign	vad_gru_input_weights_array[    1] = 32'b01000001101110000000000000000000;
	assign	vad_gru_input_weights_array[    2] = 32'b11000010111101100000000000000000;
	assign	vad_gru_input_weights_array[    3] = 32'b11000010000001000000000000000000;
	assign	vad_gru_input_weights_array[    4] = 32'b11000010101111100000000000000000;
	assign	vad_gru_input_weights_array[    5] = 32'b11000000100000000000000000000000;
	assign	vad_gru_input_weights_array[    6] = 32'b01000001000000000000000000000000;
	assign	vad_gru_input_weights_array[    7] = 32'b11000010101010000000000000000000;
	assign	vad_gru_input_weights_array[    8] = 32'b01000000100000000000000000000000;
	assign	vad_gru_input_weights_array[    9] = 32'b01000010110010100000000000000000;
	assign	vad_gru_input_weights_array[   10] = 32'b11000010111011100000000000000000;
	assign	vad_gru_input_weights_array[   11] = 32'b01000010111010000000000000000000;
	assign	vad_gru_input_weights_array[   12] = 32'b11000000100000000000000000000000;
	assign	vad_gru_input_weights_array[   13] = 32'b01000010111101100000000000000000;
	assign	vad_gru_input_weights_array[   14] = 32'b01000010110011100000000000000000;
	assign	vad_gru_input_weights_array[   15] = 32'b11000010010011000000000000000000;
	assign	vad_gru_input_weights_array[   16] = 32'b01000001111010000000000000000000;
	assign	vad_gru_input_weights_array[   17] = 32'b11000010111110000000000000000000;
	assign	vad_gru_input_weights_array[   18] = 32'b11000010111001000000000000000000;
	assign	vad_gru_input_weights_array[   19] = 32'b11000010010001000000000000000000;
	assign	vad_gru_input_weights_array[   20] = 32'b01000001111110000000000000000000;
	assign	vad_gru_input_weights_array[   21] = 32'b01000001000100000000000000000000;
	assign	vad_gru_input_weights_array[   22] = 32'b01000010100101100000000000000000;
	assign	vad_gru_input_weights_array[   23] = 32'b11000011000000000000000000000000;
	assign	vad_gru_input_weights_array[   24] = 32'b00000000000000000000000000000000;
	assign	vad_gru_input_weights_array[   25] = 32'b11000010010001000000000000000000;
	assign	vad_gru_input_weights_array[   26] = 32'b01000010000101000000000000000000;
	assign	vad_gru_input_weights_array[   27] = 32'b11000010010010000000000000000000;
	assign	vad_gru_input_weights_array[   28] = 32'b01000010001110000000000000000000;
	assign	vad_gru_input_weights_array[   29] = 32'b11000001101010000000000000000000;
	assign	vad_gru_input_weights_array[   30] = 32'b11000010011111000000000000000000;
	assign	vad_gru_input_weights_array[   31] = 32'b11000010110100000000000000000000;
	assign	vad_gru_input_weights_array[   32] = 32'b01000010010110000000000000000000;
	assign	vad_gru_input_weights_array[   33] = 32'b01000010101001000000000000000000;
	assign	vad_gru_input_weights_array[   34] = 32'b01000010000001000000000000000000;
	assign	vad_gru_input_weights_array[   35] = 32'b01000001101010000000000000000000;
	assign	vad_gru_input_weights_array[   36] = 32'b01000010100011000000000000000000;
	assign	vad_gru_input_weights_array[   37] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[   38] = 32'b11000001000100000000000000000000;
	assign	vad_gru_input_weights_array[   39] = 32'b11000010100111100000000000000000;
	assign	vad_gru_input_weights_array[   40] = 32'b11000010000111000000000000000000;
	assign	vad_gru_input_weights_array[   41] = 32'b11000001101110000000000000000000;
	assign	vad_gru_input_weights_array[   42] = 32'b11000010111111100000000000000000;
	assign	vad_gru_input_weights_array[   43] = 32'b01000010110101100000000000000000;
	assign	vad_gru_input_weights_array[   44] = 32'b01000010111101000000000000000000;
	assign	vad_gru_input_weights_array[   45] = 32'b11000010110000000000000000000000;
	assign	vad_gru_input_weights_array[   46] = 32'b11000010001110000000000000000000;
	assign	vad_gru_input_weights_array[   47] = 32'b11000001100100000000000000000000;
	assign	vad_gru_input_weights_array[   48] = 32'b11000010000111000000000000000000;
	assign	vad_gru_input_weights_array[   49] = 32'b01000001010100000000000000000000;
	assign	vad_gru_input_weights_array[   50] = 32'b11000001111000000000000000000000;
	assign	vad_gru_input_weights_array[   51] = 32'b11000010010000000000000000000000;
	assign	vad_gru_input_weights_array[   52] = 32'b01000001011000000000000000000000;
	assign	vad_gru_input_weights_array[   53] = 32'b01000010011000000000000000000000;
	assign	vad_gru_input_weights_array[   54] = 32'b11000010010100000000000000000000;
	assign	vad_gru_input_weights_array[   55] = 32'b01000010010001000000000000000000;
	assign	vad_gru_input_weights_array[   56] = 32'b10111111100000000000000000000000;
	assign	vad_gru_input_weights_array[   57] = 32'b11000010111100100000000000000000;
	assign	vad_gru_input_weights_array[   58] = 32'b01000001110010000000000000000000;
	assign	vad_gru_input_weights_array[   59] = 32'b11000001100100000000000000000000;
	assign	vad_gru_input_weights_array[   60] = 32'b11000010000100000000000000000000;
	assign	vad_gru_input_weights_array[   61] = 32'b11000010010100000000000000000000;
	assign	vad_gru_input_weights_array[   62] = 32'b11000010011001000000000000000000;
	assign	vad_gru_input_weights_array[   63] = 32'b11000001111100000000000000000000;
	assign	vad_gru_input_weights_array[   64] = 32'b01000010010110000000000000000000;
	assign	vad_gru_input_weights_array[   65] = 32'b11000010111110000000000000000000;
	assign	vad_gru_input_weights_array[   66] = 32'b11000001110100000000000000000000;
	assign	vad_gru_input_weights_array[   67] = 32'b11000010001111000000000000000000;
	assign	vad_gru_input_weights_array[   68] = 32'b01000001001000000000000000000000;
	assign	vad_gru_input_weights_array[   69] = 32'b01000010000111000000000000000000;
	assign	vad_gru_input_weights_array[   70] = 32'b01000001010000000000000000000000;
	assign	vad_gru_input_weights_array[   71] = 32'b01000000000000000000000000000000;
	assign	vad_gru_input_weights_array[   72] = 32'b01000001000100000000000000000000;
	assign	vad_gru_input_weights_array[   73] = 32'b11000010111111100000000000000000;
	assign	vad_gru_input_weights_array[   74] = 32'b11000011000000000000000000000000;
	assign	vad_gru_input_weights_array[   75] = 32'b01000010110011000000000000000000;
	assign	vad_gru_input_weights_array[   76] = 32'b01000001101010000000000000000000;
	assign	vad_gru_input_weights_array[   77] = 32'b01000001001100000000000000000000;
	assign	vad_gru_input_weights_array[   78] = 32'b11000010100000000000000000000000;
	assign	vad_gru_input_weights_array[   79] = 32'b11000010100011100000000000000000;
	assign	vad_gru_input_weights_array[   80] = 32'b01000010101100100000000000000000;
	assign	vad_gru_input_weights_array[   81] = 32'b11000010111000100000000000000000;
	assign	vad_gru_input_weights_array[   82] = 32'b11000010110111100000000000000000;
	assign	vad_gru_input_weights_array[   83] = 32'b01000010010110000000000000000000;
	assign	vad_gru_input_weights_array[   84] = 32'b01000001111110000000000000000000;
	assign	vad_gru_input_weights_array[   85] = 32'b01000010101111000000000000000000;
	assign	vad_gru_input_weights_array[   86] = 32'b01000010111100100000000000000000;
	assign	vad_gru_input_weights_array[   87] = 32'b11000010001000000000000000000000;
	assign	vad_gru_input_weights_array[   88] = 32'b01000001111100000000000000000000;
	assign	vad_gru_input_weights_array[   89] = 32'b01000010001000000000000000000000;
	assign	vad_gru_input_weights_array[   90] = 32'b11000010110110100000000000000000;
	assign	vad_gru_input_weights_array[   91] = 32'b01000010100100100000000000000000;
	assign	vad_gru_input_weights_array[   92] = 32'b11000001000100000000000000000000;
	assign	vad_gru_input_weights_array[   93] = 32'b01000010110110000000000000000000;
	assign	vad_gru_input_weights_array[   94] = 32'b11000010101110000000000000000000;
	assign	vad_gru_input_weights_array[   95] = 32'b01000000000000000000000000000000;
	assign	vad_gru_input_weights_array[   96] = 32'b11000010111111100000000000000000;
	assign	vad_gru_input_weights_array[   97] = 32'b01000010111010000000000000000000;
	assign	vad_gru_input_weights_array[   98] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[   99] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  100] = 32'b11000010111101000000000000000000;
	assign	vad_gru_input_weights_array[  101] = 32'b01000010101111100000000000000000;
	assign	vad_gru_input_weights_array[  102] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  103] = 32'b11000010000101000000000000000000;
	assign	vad_gru_input_weights_array[  104] = 32'b11000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  105] = 32'b01000001111000000000000000000000;
	assign	vad_gru_input_weights_array[  106] = 32'b01000010101100100000000000000000;
	assign	vad_gru_input_weights_array[  107] = 32'b01000001001000000000000000000000;
	assign	vad_gru_input_weights_array[  108] = 32'b01000001110000000000000000000000;
	assign	vad_gru_input_weights_array[  109] = 32'b11000010110100000000000000000000;
	assign	vad_gru_input_weights_array[  110] = 32'b11000010011110000000000000000000;
	assign	vad_gru_input_weights_array[  111] = 32'b11000010100001100000000000000000;
	assign	vad_gru_input_weights_array[  112] = 32'b11000001011000000000000000000000;
	assign	vad_gru_input_weights_array[  113] = 32'b01000010000110000000000000000000;
	assign	vad_gru_input_weights_array[  114] = 32'b01000001011000000000000000000000;
	assign	vad_gru_input_weights_array[  115] = 32'b11000010100011100000000000000000;
	assign	vad_gru_input_weights_array[  116] = 32'b01000001101100000000000000000000;
	assign	vad_gru_input_weights_array[  117] = 32'b11000010001001000000000000000000;
	assign	vad_gru_input_weights_array[  118] = 32'b01000001101000000000000000000000;
	assign	vad_gru_input_weights_array[  119] = 32'b11000010010010000000000000000000;
	assign	vad_gru_input_weights_array[  120] = 32'b01000010000111000000000000000000;
	assign	vad_gru_input_weights_array[  121] = 32'b01000010011111000000000000000000;
	assign	vad_gru_input_weights_array[  122] = 32'b01000010101011000000000000000000;
	assign	vad_gru_input_weights_array[  123] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  124] = 32'b11000001100100000000000000000000;
	assign	vad_gru_input_weights_array[  125] = 32'b01000010100111100000000000000000;
	assign	vad_gru_input_weights_array[  126] = 32'b01000000100000000000000000000000;
	assign	vad_gru_input_weights_array[  127] = 32'b11000010010011000000000000000000;
	assign	vad_gru_input_weights_array[  128] = 32'b01000000000000000000000000000000;
	assign	vad_gru_input_weights_array[  129] = 32'b01000010000001000000000000000000;
	assign	vad_gru_input_weights_array[  130] = 32'b01000010111010100000000000000000;
	assign	vad_gru_input_weights_array[  131] = 32'b11000010111000100000000000000000;
	assign	vad_gru_input_weights_array[  132] = 32'b11000010100111000000000000000000;
	assign	vad_gru_input_weights_array[  133] = 32'b01000010011000000000000000000000;
	assign	vad_gru_input_weights_array[  134] = 32'b11000010101101100000000000000000;
	assign	vad_gru_input_weights_array[  135] = 32'b01000010000101000000000000000000;
	assign	vad_gru_input_weights_array[  136] = 32'b01000010000010000000000000000000;
	assign	vad_gru_input_weights_array[  137] = 32'b11000010001101000000000000000000;
	assign	vad_gru_input_weights_array[  138] = 32'b11000010001100000000000000000000;
	assign	vad_gru_input_weights_array[  139] = 32'b11000001101100000000000000000000;
	assign	vad_gru_input_weights_array[  140] = 32'b01000001101010000000000000000000;
	assign	vad_gru_input_weights_array[  141] = 32'b11000001100000000000000000000000;
	assign	vad_gru_input_weights_array[  142] = 32'b01000010011000000000000000000000;
	assign	vad_gru_input_weights_array[  143] = 32'b01000001111100000000000000000000;
	assign	vad_gru_input_weights_array[  144] = 32'b11000010101010000000000000000000;
	assign	vad_gru_input_weights_array[  145] = 32'b11000010100111100000000000000000;
	assign	vad_gru_input_weights_array[  146] = 32'b01000010000110000000000000000000;
	assign	vad_gru_input_weights_array[  147] = 32'b11000010100101000000000000000000;
	assign	vad_gru_input_weights_array[  148] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  149] = 32'b01000001000100000000000000000000;
	assign	vad_gru_input_weights_array[  150] = 32'b11000001110010000000000000000000;
	assign	vad_gru_input_weights_array[  151] = 32'b01000000000000000000000000000000;
	assign	vad_gru_input_weights_array[  152] = 32'b01000010101001000000000000000000;
	assign	vad_gru_input_weights_array[  153] = 32'b01000010011101000000000000000000;
	assign	vad_gru_input_weights_array[  154] = 32'b01000001110010000000000000000000;
	assign	vad_gru_input_weights_array[  155] = 32'b11000001110100000000000000000000;
	assign	vad_gru_input_weights_array[  156] = 32'b01000001110100000000000000000000;
	assign	vad_gru_input_weights_array[  157] = 32'b01000001001100000000000000000000;
	assign	vad_gru_input_weights_array[  158] = 32'b01000010111010100000000000000000;
	assign	vad_gru_input_weights_array[  159] = 32'b11000010100000100000000000000000;
	assign	vad_gru_input_weights_array[  160] = 32'b01000001010000000000000000000000;
	assign	vad_gru_input_weights_array[  161] = 32'b11000010011010000000000000000000;
	assign	vad_gru_input_weights_array[  162] = 32'b01000010001010000000000000000000;
	assign	vad_gru_input_weights_array[  163] = 32'b11000010011110000000000000000000;
	assign	vad_gru_input_weights_array[  164] = 32'b11000010101110100000000000000000;
	assign	vad_gru_input_weights_array[  165] = 32'b01000001001100000000000000000000;
	assign	vad_gru_input_weights_array[  166] = 32'b01000001001100000000000000000000;
	assign	vad_gru_input_weights_array[  167] = 32'b01000010111110000000000000000000;
	assign	vad_gru_input_weights_array[  168] = 32'b11000010111101100000000000000000;
	assign	vad_gru_input_weights_array[  169] = 32'b01000010101000000000000000000000;
	assign	vad_gru_input_weights_array[  170] = 32'b11000010111110100000000000000000;
	assign	vad_gru_input_weights_array[  171] = 32'b01000001001100000000000000000000;
	assign	vad_gru_input_weights_array[  172] = 32'b11000010101101000000000000000000;
	assign	vad_gru_input_weights_array[  173] = 32'b01000010001010000000000000000000;
	assign	vad_gru_input_weights_array[  174] = 32'b01000010101111000000000000000000;
	assign	vad_gru_input_weights_array[  175] = 32'b01000000100000000000000000000000;
	assign	vad_gru_input_weights_array[  176] = 32'b11000010110110100000000000000000;
	assign	vad_gru_input_weights_array[  177] = 32'b10111111100000000000000000000000;
	assign	vad_gru_input_weights_array[  178] = 32'b01000010101010100000000000000000;
	assign	vad_gru_input_weights_array[  179] = 32'b11000010010100000000000000000000;
	assign	vad_gru_input_weights_array[  180] = 32'b01000010001101000000000000000000;
	assign	vad_gru_input_weights_array[  181] = 32'b11000001110100000000000000000000;
	assign	vad_gru_input_weights_array[  182] = 32'b11000001110110000000000000000000;
	assign	vad_gru_input_weights_array[  183] = 32'b01000010100110100000000000000000;
	assign	vad_gru_input_weights_array[  184] = 32'b11000000101000000000000000000000;
	assign	vad_gru_input_weights_array[  185] = 32'b01000001111100000000000000000000;
	assign	vad_gru_input_weights_array[  186] = 32'b01000010101101000000000000000000;
	assign	vad_gru_input_weights_array[  187] = 32'b00000000000000000000000000000000;
	assign	vad_gru_input_weights_array[  188] = 32'b01000010101111100000000000000000;
	assign	vad_gru_input_weights_array[  189] = 32'b11000000111000000000000000000000;
	assign	vad_gru_input_weights_array[  190] = 32'b01000010010101000000000000000000;
	assign	vad_gru_input_weights_array[  191] = 32'b01000001111010000000000000000000;
	assign	vad_gru_input_weights_array[  192] = 32'b11000010101001000000000000000000;
	assign	vad_gru_input_weights_array[  193] = 32'b01000001101100000000000000000000;
	assign	vad_gru_input_weights_array[  194] = 32'b11000001000100000000000000000000;
	assign	vad_gru_input_weights_array[  195] = 32'b01000010100101000000000000000000;
	assign	vad_gru_input_weights_array[  196] = 32'b01000000000000000000000000000000;
	assign	vad_gru_input_weights_array[  197] = 32'b11000001010000000000000000000000;
	assign	vad_gru_input_weights_array[  198] = 32'b11000010100100100000000000000000;
	assign	vad_gru_input_weights_array[  199] = 32'b01000010111001000000000000000000;
	assign	vad_gru_input_weights_array[  200] = 32'b01000010110000100000000000000000;
	assign	vad_gru_input_weights_array[  201] = 32'b11000010100000000000000000000000;
	assign	vad_gru_input_weights_array[  202] = 32'b01000010111101000000000000000000;
	assign	vad_gru_input_weights_array[  203] = 32'b11000010100110100000000000000000;
	assign	vad_gru_input_weights_array[  204] = 32'b01000010001011000000000000000000;
	assign	vad_gru_input_weights_array[  205] = 32'b01000010101101100000000000000000;
	assign	vad_gru_input_weights_array[  206] = 32'b01000010101011000000000000000000;
	assign	vad_gru_input_weights_array[  207] = 32'b01000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  208] = 32'b01000010110101000000000000000000;
	assign	vad_gru_input_weights_array[  209] = 32'b01000010100100000000000000000000;
	assign	vad_gru_input_weights_array[  210] = 32'b01000010101101000000000000000000;
	assign	vad_gru_input_weights_array[  211] = 32'b11000010001011000000000000000000;
	assign	vad_gru_input_weights_array[  212] = 32'b01000010001110000000000000000000;
	assign	vad_gru_input_weights_array[  213] = 32'b01000010110000000000000000000000;
	assign	vad_gru_input_weights_array[  214] = 32'b11000010010011000000000000000000;
	assign	vad_gru_input_weights_array[  215] = 32'b01000001101010000000000000000000;
	assign	vad_gru_input_weights_array[  216] = 32'b01000001101100000000000000000000;
	assign	vad_gru_input_weights_array[  217] = 32'b01000010100010000000000000000000;
	assign	vad_gru_input_weights_array[  218] = 32'b01000001101100000000000000000000;
	assign	vad_gru_input_weights_array[  219] = 32'b01000010001001000000000000000000;
	assign	vad_gru_input_weights_array[  220] = 32'b01000010100111100000000000000000;
	assign	vad_gru_input_weights_array[  221] = 32'b01000010100101100000000000000000;
	assign	vad_gru_input_weights_array[  222] = 32'b11000010001110000000000000000000;
	assign	vad_gru_input_weights_array[  223] = 32'b11000010110100100000000000000000;
	assign	vad_gru_input_weights_array[  224] = 32'b01000001101110000000000000000000;
	assign	vad_gru_input_weights_array[  225] = 32'b11000010111010000000000000000000;
	assign	vad_gru_input_weights_array[  226] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  227] = 32'b11000010111101100000000000000000;
	assign	vad_gru_input_weights_array[  228] = 32'b01000010110011000000000000000000;
	assign	vad_gru_input_weights_array[  229] = 32'b01000010011001000000000000000000;
	assign	vad_gru_input_weights_array[  230] = 32'b01000010101010100000000000000000;
	assign	vad_gru_input_weights_array[  231] = 32'b01000001001000000000000000000000;
	assign	vad_gru_input_weights_array[  232] = 32'b11000001111010000000000000000000;
	assign	vad_gru_input_weights_array[  233] = 32'b01000010000010000000000000000000;
	assign	vad_gru_input_weights_array[  234] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[  235] = 32'b01000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  236] = 32'b01000010111110000000000000000000;
	assign	vad_gru_input_weights_array[  237] = 32'b01000010101000100000000000000000;
	assign	vad_gru_input_weights_array[  238] = 32'b11000001011100000000000000000000;
	assign	vad_gru_input_weights_array[  239] = 32'b01000010010110000000000000000000;
	assign	vad_gru_input_weights_array[  240] = 32'b01000010110000000000000000000000;
	assign	vad_gru_input_weights_array[  241] = 32'b11000011000000000000000000000000;
	assign	vad_gru_input_weights_array[  242] = 32'b01000010000111000000000000000000;
	assign	vad_gru_input_weights_array[  243] = 32'b11000010111110000000000000000000;
	assign	vad_gru_input_weights_array[  244] = 32'b01000010110011100000000000000000;
	assign	vad_gru_input_weights_array[  245] = 32'b01000010100101000000000000000000;
	assign	vad_gru_input_weights_array[  246] = 32'b01000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  247] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  248] = 32'b11000010010010000000000000000000;
	assign	vad_gru_input_weights_array[  249] = 32'b11000010100011100000000000000000;
	assign	vad_gru_input_weights_array[  250] = 32'b11000010111101000000000000000000;
	assign	vad_gru_input_weights_array[  251] = 32'b11000010100000000000000000000000;
	assign	vad_gru_input_weights_array[  252] = 32'b01000010101110100000000000000000;
	assign	vad_gru_input_weights_array[  253] = 32'b11000010100101100000000000000000;
	assign	vad_gru_input_weights_array[  254] = 32'b01000010100011100000000000000000;
	assign	vad_gru_input_weights_array[  255] = 32'b01000010110100100000000000000000;
	assign	vad_gru_input_weights_array[  256] = 32'b01000010111101000000000000000000;
	assign	vad_gru_input_weights_array[  257] = 32'b01000010111101100000000000000000;
	assign	vad_gru_input_weights_array[  258] = 32'b01000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  259] = 32'b01000010111101000000000000000000;
	assign	vad_gru_input_weights_array[  260] = 32'b11000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  261] = 32'b01000010000001000000000000000000;
	assign	vad_gru_input_weights_array[  262] = 32'b11000010011111000000000000000000;
	assign	vad_gru_input_weights_array[  263] = 32'b11000010100101000000000000000000;
	assign	vad_gru_input_weights_array[  264] = 32'b01000010111110000000000000000000;
	assign	vad_gru_input_weights_array[  265] = 32'b11000010100011100000000000000000;
	assign	vad_gru_input_weights_array[  266] = 32'b01000010000001000000000000000000;
	assign	vad_gru_input_weights_array[  267] = 32'b01000010001001000000000000000000;
	assign	vad_gru_input_weights_array[  268] = 32'b11000010011000000000000000000000;
	assign	vad_gru_input_weights_array[  269] = 32'b01000001100110000000000000000000;
	assign	vad_gru_input_weights_array[  270] = 32'b01000000110000000000000000000000;
	assign	vad_gru_input_weights_array[  271] = 32'b01000010100000100000000000000000;
	assign	vad_gru_input_weights_array[  272] = 32'b01000010001001000000000000000000;
	assign	vad_gru_input_weights_array[  273] = 32'b01000010101101000000000000000000;
	assign	vad_gru_input_weights_array[  274] = 32'b11000010111010000000000000000000;
	assign	vad_gru_input_weights_array[  275] = 32'b11000000010000000000000000000000;
	assign	vad_gru_input_weights_array[  276] = 32'b11000010001110000000000000000000;
	assign	vad_gru_input_weights_array[  277] = 32'b01000010100101100000000000000000;
	assign	vad_gru_input_weights_array[  278] = 32'b11000001010100000000000000000000;
	assign	vad_gru_input_weights_array[  279] = 32'b01000010110001000000000000000000;
	assign	vad_gru_input_weights_array[  280] = 32'b11000010100101000000000000000000;
	assign	vad_gru_input_weights_array[  281] = 32'b11000010001010000000000000000000;
	assign	vad_gru_input_weights_array[  282] = 32'b01000010100101000000000000000000;
	assign	vad_gru_input_weights_array[  283] = 32'b11000010101111100000000000000000;
	assign	vad_gru_input_weights_array[  284] = 32'b11000010110000000000000000000000;
	assign	vad_gru_input_weights_array[  285] = 32'b01000010101000100000000000000000;
	assign	vad_gru_input_weights_array[  286] = 32'b01000001110000000000000000000000;
	assign	vad_gru_input_weights_array[  287] = 32'b01000010000000000000000000000000;
	assign	vad_gru_input_weights_array[  288] = 32'b11000001100110000000000000000000;
	assign	vad_gru_input_weights_array[  289] = 32'b11000010111101100000000000000000;
	assign	vad_gru_input_weights_array[  290] = 32'b01000010100101000000000000000000;
	assign	vad_gru_input_weights_array[  291] = 32'b01000010010111000000000000000000;
	assign	vad_gru_input_weights_array[  292] = 32'b01000010110110100000000000000000;
	assign	vad_gru_input_weights_array[  293] = 32'b01000010111001100000000000000000;
	assign	vad_gru_input_weights_array[  294] = 32'b00000000000000000000000000000000;
	assign	vad_gru_input_weights_array[  295] = 32'b01000010000000000000000000000000;
	assign	vad_gru_input_weights_array[  296] = 32'b01000010000001000000000000000000;
	assign	vad_gru_input_weights_array[  297] = 32'b01000001010000000000000000000000;
	assign	vad_gru_input_weights_array[  298] = 32'b11000001101000000000000000000000;
	assign	vad_gru_input_weights_array[  299] = 32'b01000001000100000000000000000000;
	assign	vad_gru_input_weights_array[  300] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  301] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  302] = 32'b11000010011101000000000000000000;
	assign	vad_gru_input_weights_array[  303] = 32'b01000010100111100000000000000000;
	assign	vad_gru_input_weights_array[  304] = 32'b11000010010000000000000000000000;
	assign	vad_gru_input_weights_array[  305] = 32'b11000010010110000000000000000000;
	assign	vad_gru_input_weights_array[  306] = 32'b11000010010001000000000000000000;
	assign	vad_gru_input_weights_array[  307] = 32'b01000010110010100000000000000000;
	assign	vad_gru_input_weights_array[  308] = 32'b11000001000100000000000000000000;
	assign	vad_gru_input_weights_array[  309] = 32'b01000001110110000000000000000000;
	assign	vad_gru_input_weights_array[  310] = 32'b11000010110101000000000000000000;
	assign	vad_gru_input_weights_array[  311] = 32'b01000010100101000000000000000000;
	assign	vad_gru_input_weights_array[  312] = 32'b01000010111011100000000000000000;
	assign	vad_gru_input_weights_array[  313] = 32'b01000010100110100000000000000000;
	assign	vad_gru_input_weights_array[  314] = 32'b01000010101011100000000000000000;
	assign	vad_gru_input_weights_array[  315] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  316] = 32'b11000001110000000000000000000000;
	assign	vad_gru_input_weights_array[  317] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  318] = 32'b01000010111110000000000000000000;
	assign	vad_gru_input_weights_array[  319] = 32'b01000001111110000000000000000000;
	assign	vad_gru_input_weights_array[  320] = 32'b01000010000010000000000000000000;
	assign	vad_gru_input_weights_array[  321] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  322] = 32'b01000010001000000000000000000000;
	assign	vad_gru_input_weights_array[  323] = 32'b01000000010000000000000000000000;
	assign	vad_gru_input_weights_array[  324] = 32'b11000010101101000000000000000000;
	assign	vad_gru_input_weights_array[  325] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  326] = 32'b01000001101110000000000000000000;
	assign	vad_gru_input_weights_array[  327] = 32'b01000010011001000000000000000000;
	assign	vad_gru_input_weights_array[  328] = 32'b11000010010101000000000000000000;
	assign	vad_gru_input_weights_array[  329] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  330] = 32'b11000010100010100000000000000000;
	assign	vad_gru_input_weights_array[  331] = 32'b11000010101100000000000000000000;
	assign	vad_gru_input_weights_array[  332] = 32'b11000010000001000000000000000000;
	assign	vad_gru_input_weights_array[  333] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  334] = 32'b01000001100110000000000000000000;
	assign	vad_gru_input_weights_array[  335] = 32'b11000010001110000000000000000000;
	assign	vad_gru_input_weights_array[  336] = 32'b11000001000100000000000000000000;
	assign	vad_gru_input_weights_array[  337] = 32'b11000010111110100000000000000000;
	assign	vad_gru_input_weights_array[  338] = 32'b01000001010100000000000000000000;
	assign	vad_gru_input_weights_array[  339] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  340] = 32'b11000010111000100000000000000000;
	assign	vad_gru_input_weights_array[  341] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  342] = 32'b11000010001001000000000000000000;
	assign	vad_gru_input_weights_array[  343] = 32'b01000010001110000000000000000000;
	assign	vad_gru_input_weights_array[  344] = 32'b01000010110101000000000000000000;
	assign	vad_gru_input_weights_array[  345] = 32'b11000010011110000000000000000000;
	assign	vad_gru_input_weights_array[  346] = 32'b01000000010000000000000000000000;
	assign	vad_gru_input_weights_array[  347] = 32'b11000001001000000000000000000000;
	assign	vad_gru_input_weights_array[  348] = 32'b01000010110111100000000000000000;
	assign	vad_gru_input_weights_array[  349] = 32'b01000010010001000000000000000000;
	assign	vad_gru_input_weights_array[  350] = 32'b11000010000010000000000000000000;
	assign	vad_gru_input_weights_array[  351] = 32'b11000001110000000000000000000000;
	assign	vad_gru_input_weights_array[  352] = 32'b11000001101000000000000000000000;
	assign	vad_gru_input_weights_array[  353] = 32'b11000010111000000000000000000000;
	assign	vad_gru_input_weights_array[  354] = 32'b01000001001100000000000000000000;
	assign	vad_gru_input_weights_array[  355] = 32'b01000010110010100000000000000000;
	assign	vad_gru_input_weights_array[  356] = 32'b11000010010010000000000000000000;
	assign	vad_gru_input_weights_array[  357] = 32'b11000010000010000000000000000000;
	assign	vad_gru_input_weights_array[  358] = 32'b01000010010010000000000000000000;
	assign	vad_gru_input_weights_array[  359] = 32'b01000010100000100000000000000000;
	assign	vad_gru_input_weights_array[  360] = 32'b11000010100000000000000000000000;
	assign	vad_gru_input_weights_array[  361] = 32'b11000010110101000000000000000000;
	assign	vad_gru_input_weights_array[  362] = 32'b01000010100011000000000000000000;
	assign	vad_gru_input_weights_array[  363] = 32'b11000010010000000000000000000000;
	assign	vad_gru_input_weights_array[  364] = 32'b01000010011100000000000000000000;
	assign	vad_gru_input_weights_array[  365] = 32'b01000001000100000000000000000000;
	assign	vad_gru_input_weights_array[  366] = 32'b11000010111101000000000000000000;
	assign	vad_gru_input_weights_array[  367] = 32'b11000010001101000000000000000000;
	assign	vad_gru_input_weights_array[  368] = 32'b01000001011100000000000000000000;
	assign	vad_gru_input_weights_array[  369] = 32'b11000010111000000000000000000000;
	assign	vad_gru_input_weights_array[  370] = 32'b11000001110100000000000000000000;
	assign	vad_gru_input_weights_array[  371] = 32'b11000000100000000000000000000000;
	assign	vad_gru_input_weights_array[  372] = 32'b00111111100000000000000000000000;
	assign	vad_gru_input_weights_array[  373] = 32'b01000010000111000000000000000000;
	assign	vad_gru_input_weights_array[  374] = 32'b01000001101110000000000000000000;
	assign	vad_gru_input_weights_array[  375] = 32'b01000010011010000000000000000000;
	assign	vad_gru_input_weights_array[  376] = 32'b11000010001101000000000000000000;
	assign	vad_gru_input_weights_array[  377] = 32'b11000010101000000000000000000000;
	assign	vad_gru_input_weights_array[  378] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  379] = 32'b01000010101001000000000000000000;
	assign	vad_gru_input_weights_array[  380] = 32'b01000010011010000000000000000000;
	assign	vad_gru_input_weights_array[  381] = 32'b01000001111100000000000000000000;
	assign	vad_gru_input_weights_array[  382] = 32'b11000010101111000000000000000000;
	assign	vad_gru_input_weights_array[  383] = 32'b11000010111011100000000000000000;
	assign	vad_gru_input_weights_array[  384] = 32'b01000010010011000000000000000000;
	assign	vad_gru_input_weights_array[  385] = 32'b11000010101100100000000000000000;
	assign	vad_gru_input_weights_array[  386] = 32'b01000010101111100000000000000000;
	assign	vad_gru_input_weights_array[  387] = 32'b11000010110101100000000000000000;
	assign	vad_gru_input_weights_array[  388] = 32'b01000001111100000000000000000000;
	assign	vad_gru_input_weights_array[  389] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  390] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[  391] = 32'b01000010011010000000000000000000;
	assign	vad_gru_input_weights_array[  392] = 32'b11000010010100000000000000000000;
	assign	vad_gru_input_weights_array[  393] = 32'b11000010001010000000000000000000;
	assign	vad_gru_input_weights_array[  394] = 32'b11000010000110000000000000000000;
	assign	vad_gru_input_weights_array[  395] = 32'b11000001101000000000000000000000;
	assign	vad_gru_input_weights_array[  396] = 32'b11000010111101000000000000000000;
	assign	vad_gru_input_weights_array[  397] = 32'b01000010111001100000000000000000;
	assign	vad_gru_input_weights_array[  398] = 32'b01000010000111000000000000000000;
	assign	vad_gru_input_weights_array[  399] = 32'b11000001110100000000000000000000;
	assign	vad_gru_input_weights_array[  400] = 32'b01000000101000000000000000000000;
	assign	vad_gru_input_weights_array[  401] = 32'b01000010100100100000000000000000;
	assign	vad_gru_input_weights_array[  402] = 32'b01000001010100000000000000000000;
	assign	vad_gru_input_weights_array[  403] = 32'b11000010000111000000000000000000;
	assign	vad_gru_input_weights_array[  404] = 32'b01000010001011000000000000000000;
	assign	vad_gru_input_weights_array[  405] = 32'b11000001101110000000000000000000;
	assign	vad_gru_input_weights_array[  406] = 32'b11000001101000000000000000000000;
	assign	vad_gru_input_weights_array[  407] = 32'b11000010111110100000000000000000;
	assign	vad_gru_input_weights_array[  408] = 32'b01000001101110000000000000000000;
	assign	vad_gru_input_weights_array[  409] = 32'b01000010000011000000000000000000;
	assign	vad_gru_input_weights_array[  410] = 32'b01000010010101000000000000000000;
	assign	vad_gru_input_weights_array[  411] = 32'b11000010011101000000000000000000;
	assign	vad_gru_input_weights_array[  412] = 32'b11000010100001000000000000000000;
	assign	vad_gru_input_weights_array[  413] = 32'b01000010100100000000000000000000;
	assign	vad_gru_input_weights_array[  414] = 32'b11000001101000000000000000000000;
	assign	vad_gru_input_weights_array[  415] = 32'b01000010000001000000000000000000;
	assign	vad_gru_input_weights_array[  416] = 32'b01000001000000000000000000000000;
	assign	vad_gru_input_weights_array[  417] = 32'b01000010000011000000000000000000;
	assign	vad_gru_input_weights_array[  418] = 32'b01000000100000000000000000000000;
	assign	vad_gru_input_weights_array[  419] = 32'b01000000111000000000000000000000;
	assign	vad_gru_input_weights_array[  420] = 32'b01000001100100000000000000000000;
	assign	vad_gru_input_weights_array[  421] = 32'b01000001100110000000000000000000;
	assign	vad_gru_input_weights_array[  422] = 32'b01000001100000000000000000000000;
	assign	vad_gru_input_weights_array[  423] = 32'b11000010001101000000000000000000;
	assign	vad_gru_input_weights_array[  424] = 32'b11000010010010000000000000000000;
	assign	vad_gru_input_weights_array[  425] = 32'b11000010100011100000000000000000;
	assign	vad_gru_input_weights_array[  426] = 32'b01000001111110000000000000000000;
	assign	vad_gru_input_weights_array[  427] = 32'b11000001111010000000000000000000;
	assign	vad_gru_input_weights_array[  428] = 32'b11000010001001000000000000000000;
	assign	vad_gru_input_weights_array[  429] = 32'b11000001110110000000000000000000;
	assign	vad_gru_input_weights_array[  430] = 32'b01000001001000000000000000000000;
	assign	vad_gru_input_weights_array[  431] = 32'b01000001011000000000000000000000;
	assign	vad_gru_input_weights_array[  432] = 32'b01000001110110000000000000000000;
	assign	vad_gru_input_weights_array[  433] = 32'b01000001000100000000000000000000;
	assign	vad_gru_input_weights_array[  434] = 32'b11000001101110000000000000000000;
	assign	vad_gru_input_weights_array[  435] = 32'b01000010110001000000000000000000;
	assign	vad_gru_input_weights_array[  436] = 32'b01000000110000000000000000000000;
	assign	vad_gru_input_weights_array[  437] = 32'b11000010101111000000000000000000;
	assign	vad_gru_input_weights_array[  438] = 32'b01000010101110000000000000000000;
	assign	vad_gru_input_weights_array[  439] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  440] = 32'b11000010111001000000000000000000;
	assign	vad_gru_input_weights_array[  441] = 32'b01000010011011000000000000000000;
	assign	vad_gru_input_weights_array[  442] = 32'b11000001110100000000000000000000;
	assign	vad_gru_input_weights_array[  443] = 32'b11000010110010000000000000000000;
	assign	vad_gru_input_weights_array[  444] = 32'b11000010011110000000000000000000;
	assign	vad_gru_input_weights_array[  445] = 32'b11000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  446] = 32'b11000001100010000000000000000000;
	assign	vad_gru_input_weights_array[  447] = 32'b11000010101010100000000000000000;
	assign	vad_gru_input_weights_array[  448] = 32'b11000010011100000000000000000000;
	assign	vad_gru_input_weights_array[  449] = 32'b01000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  450] = 32'b11000010001010000000000000000000;
	assign	vad_gru_input_weights_array[  451] = 32'b11000000110000000000000000000000;
	assign	vad_gru_input_weights_array[  452] = 32'b01000010000001000000000000000000;
	assign	vad_gru_input_weights_array[  453] = 32'b11000010111100000000000000000000;
	assign	vad_gru_input_weights_array[  454] = 32'b11000001110100000000000000000000;
	assign	vad_gru_input_weights_array[  455] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  456] = 32'b11000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  457] = 32'b11000010000011000000000000000000;
	assign	vad_gru_input_weights_array[  458] = 32'b11000010111001000000000000000000;
	assign	vad_gru_input_weights_array[  459] = 32'b11000001111110000000000000000000;
	assign	vad_gru_input_weights_array[  460] = 32'b01000001110010000000000000000000;
	assign	vad_gru_input_weights_array[  461] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  462] = 32'b11000010110010000000000000000000;
	assign	vad_gru_input_weights_array[  463] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  464] = 32'b11000010100000000000000000000000;
	assign	vad_gru_input_weights_array[  465] = 32'b11000010001110000000000000000000;
	assign	vad_gru_input_weights_array[  466] = 32'b11000001111110000000000000000000;
	assign	vad_gru_input_weights_array[  467] = 32'b01000001111100000000000000000000;
	assign	vad_gru_input_weights_array[  468] = 32'b01000001110010000000000000000000;
	assign	vad_gru_input_weights_array[  469] = 32'b11000010100101000000000000000000;
	assign	vad_gru_input_weights_array[  470] = 32'b11000010110111100000000000000000;
	assign	vad_gru_input_weights_array[  471] = 32'b11000010110000100000000000000000;
	assign	vad_gru_input_weights_array[  472] = 32'b11000010101000100000000000000000;
	assign	vad_gru_input_weights_array[  473] = 32'b11000010110100000000000000000000;
	assign	vad_gru_input_weights_array[  474] = 32'b11000010111001000000000000000000;
	assign	vad_gru_input_weights_array[  475] = 32'b11000001100110000000000000000000;
	assign	vad_gru_input_weights_array[  476] = 32'b11000001000100000000000000000000;
	assign	vad_gru_input_weights_array[  477] = 32'b11000010111010000000000000000000;
	assign	vad_gru_input_weights_array[  478] = 32'b11000010100010100000000000000000;
	assign	vad_gru_input_weights_array[  479] = 32'b01000001101100000000000000000000;
	assign	vad_gru_input_weights_array[  480] = 32'b01000001111100000000000000000000;
	assign	vad_gru_input_weights_array[  481] = 32'b01000010011011000000000000000000;
	assign	vad_gru_input_weights_array[  482] = 32'b01000001000000000000000000000000;
	assign	vad_gru_input_weights_array[  483] = 32'b11000010010011000000000000000000;
	assign	vad_gru_input_weights_array[  484] = 32'b01000001100000000000000000000000;
	assign	vad_gru_input_weights_array[  485] = 32'b11000010110000100000000000000000;
	assign	vad_gru_input_weights_array[  486] = 32'b01000001100100000000000000000000;
	assign	vad_gru_input_weights_array[  487] = 32'b11000000100000000000000000000000;
	assign	vad_gru_input_weights_array[  488] = 32'b11000010101100100000000000000000;
	assign	vad_gru_input_weights_array[  489] = 32'b01000010101000000000000000000000;
	assign	vad_gru_input_weights_array[  490] = 32'b11000010010010000000000000000000;
	assign	vad_gru_input_weights_array[  491] = 32'b01000000010000000000000000000000;
	assign	vad_gru_input_weights_array[  492] = 32'b01000010000100000000000000000000;
	assign	vad_gru_input_weights_array[  493] = 32'b11000010100001100000000000000000;
	assign	vad_gru_input_weights_array[  494] = 32'b01000010011000000000000000000000;
	assign	vad_gru_input_weights_array[  495] = 32'b01000010100010100000000000000000;
	assign	vad_gru_input_weights_array[  496] = 32'b11000001110100000000000000000000;
	assign	vad_gru_input_weights_array[  497] = 32'b01000010110101100000000000000000;
	assign	vad_gru_input_weights_array[  498] = 32'b11000001001000000000000000000000;
	assign	vad_gru_input_weights_array[  499] = 32'b01000010011010000000000000000000;
	assign	vad_gru_input_weights_array[  500] = 32'b11000001111000000000000000000000;
	assign	vad_gru_input_weights_array[  501] = 32'b11000000100000000000000000000000;
	assign	vad_gru_input_weights_array[  502] = 32'b11000010011001000000000000000000;
	assign	vad_gru_input_weights_array[  503] = 32'b11000010100100000000000000000000;
	assign	vad_gru_input_weights_array[  504] = 32'b11000010110111100000000000000000;
	assign	vad_gru_input_weights_array[  505] = 32'b00000000000000000000000000000000;
	assign	vad_gru_input_weights_array[  506] = 32'b11000010100101100000000000000000;
	assign	vad_gru_input_weights_array[  507] = 32'b11000010111011100000000000000000;
	assign	vad_gru_input_weights_array[  508] = 32'b01000001011000000000000000000000;
	assign	vad_gru_input_weights_array[  509] = 32'b11000010100101100000000000000000;
	assign	vad_gru_input_weights_array[  510] = 32'b11000010010001000000000000000000;
	assign	vad_gru_input_weights_array[  511] = 32'b11000010100001000000000000000000;
	assign	vad_gru_input_weights_array[  512] = 32'b11000010010001000000000000000000;
	assign	vad_gru_input_weights_array[  513] = 32'b01000001000000000000000000000000;
	assign	vad_gru_input_weights_array[  514] = 32'b11000010111100100000000000000000;
	assign	vad_gru_input_weights_array[  515] = 32'b01000001101100000000000000000000;
	assign	vad_gru_input_weights_array[  516] = 32'b11000010010110000000000000000000;
	assign	vad_gru_input_weights_array[  517] = 32'b01000010111100100000000000000000;
	assign	vad_gru_input_weights_array[  518] = 32'b01000001111100000000000000000000;
	assign	vad_gru_input_weights_array[  519] = 32'b01000010010110000000000000000000;
	assign	vad_gru_input_weights_array[  520] = 32'b11000001110100000000000000000000;
	assign	vad_gru_input_weights_array[  521] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  522] = 32'b11000010111101100000000000000000;
	assign	vad_gru_input_weights_array[  523] = 32'b01000010011000000000000000000000;
	assign	vad_gru_input_weights_array[  524] = 32'b01000000101000000000000000000000;
	assign	vad_gru_input_weights_array[  525] = 32'b01000010010000000000000000000000;
	assign	vad_gru_input_weights_array[  526] = 32'b01000001101010000000000000000000;
	assign	vad_gru_input_weights_array[  527] = 32'b11000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  528] = 32'b11000001001100000000000000000000;
	assign	vad_gru_input_weights_array[  529] = 32'b01000001101110000000000000000000;
	assign	vad_gru_input_weights_array[  530] = 32'b01000001110010000000000000000000;
	assign	vad_gru_input_weights_array[  531] = 32'b11000010101001000000000000000000;
	assign	vad_gru_input_weights_array[  532] = 32'b01000000110000000000000000000000;
	assign	vad_gru_input_weights_array[  533] = 32'b11000001110010000000000000000000;
	assign	vad_gru_input_weights_array[  534] = 32'b01000010111011100000000000000000;
	assign	vad_gru_input_weights_array[  535] = 32'b01000010100111000000000000000000;
	assign	vad_gru_input_weights_array[  536] = 32'b01000000100000000000000000000000;
	assign	vad_gru_input_weights_array[  537] = 32'b11000010110100000000000000000000;
	assign	vad_gru_input_weights_array[  538] = 32'b01000001110110000000000000000000;
	assign	vad_gru_input_weights_array[  539] = 32'b01000010011101000000000000000000;
	assign	vad_gru_input_weights_array[  540] = 32'b11000010010000000000000000000000;
	assign	vad_gru_input_weights_array[  541] = 32'b01000010000101000000000000000000;
	assign	vad_gru_input_weights_array[  542] = 32'b11000001010100000000000000000000;
	assign	vad_gru_input_weights_array[  543] = 32'b11000010010100000000000000000000;
	assign	vad_gru_input_weights_array[  544] = 32'b01000010010010000000000000000000;
	assign	vad_gru_input_weights_array[  545] = 32'b11000010010010000000000000000000;
	assign	vad_gru_input_weights_array[  546] = 32'b01000010001100000000000000000000;
	assign	vad_gru_input_weights_array[  547] = 32'b10111111100000000000000000000000;
	assign	vad_gru_input_weights_array[  548] = 32'b11000001101100000000000000000000;
	assign	vad_gru_input_weights_array[  549] = 32'b11000010001011000000000000000000;
	assign	vad_gru_input_weights_array[  550] = 32'b11000010011011000000000000000000;
	assign	vad_gru_input_weights_array[  551] = 32'b11000010100111000000000000000000;
	assign	vad_gru_input_weights_array[  552] = 32'b11000010100001100000000000000000;
	assign	vad_gru_input_weights_array[  553] = 32'b11000010000000000000000000000000;
	assign	vad_gru_input_weights_array[  554] = 32'b11000001110100000000000000000000;
	assign	vad_gru_input_weights_array[  555] = 32'b01000001000100000000000000000000;
	assign	vad_gru_input_weights_array[  556] = 32'b11000000010000000000000000000000;
	assign	vad_gru_input_weights_array[  557] = 32'b01000010001000000000000000000000;
	assign	vad_gru_input_weights_array[  558] = 32'b01000001100000000000000000000000;
	assign	vad_gru_input_weights_array[  559] = 32'b01000001100110000000000000000000;
	assign	vad_gru_input_weights_array[  560] = 32'b01000000010000000000000000000000;
	assign	vad_gru_input_weights_array[  561] = 32'b11000001000100000000000000000000;
	assign	vad_gru_input_weights_array[  562] = 32'b01000001101000000000000000000000;
	assign	vad_gru_input_weights_array[  563] = 32'b11000000110000000000000000000000;
	assign	vad_gru_input_weights_array[  564] = 32'b11000010000101000000000000000000;
	assign	vad_gru_input_weights_array[  565] = 32'b01000001111000000000000000000000;
	assign	vad_gru_input_weights_array[  566] = 32'b01000010000111000000000000000000;
	assign	vad_gru_input_weights_array[  567] = 32'b01000001100010000000000000000000;
	assign	vad_gru_input_weights_array[  568] = 32'b11000001100110000000000000000000;
	assign	vad_gru_input_weights_array[  569] = 32'b11000001001000000000000000000000;
	assign	vad_gru_input_weights_array[  570] = 32'b00111111100000000000000000000000;
	assign	vad_gru_input_weights_array[  571] = 32'b01000000110000000000000000000000;
	assign	vad_gru_input_weights_array[  572] = 32'b11000010011011000000000000000000;
	assign	vad_gru_input_weights_array[  573] = 32'b01000010100101000000000000000000;
	assign	vad_gru_input_weights_array[  574] = 32'b01000010001111000000000000000000;
	assign	vad_gru_input_weights_array[  575] = 32'b01000000010000000000000000000000;
	assign	vad_gru_input_weights_array[  576] = 32'b11000010111011100000000000000000;
	assign	vad_gru_input_weights_array[  577] = 32'b00000000000000000000000000000000;
	assign	vad_gru_input_weights_array[  578] = 32'b11000011000000000000000000000000;
	assign	vad_gru_input_weights_array[  579] = 32'b11000010110101100000000000000000;
	assign	vad_gru_input_weights_array[  580] = 32'b11000001110010000000000000000000;
	assign	vad_gru_input_weights_array[  581] = 32'b11000001101100000000000000000000;
	assign	vad_gru_input_weights_array[  582] = 32'b11000010100010100000000000000000;
	assign	vad_gru_input_weights_array[  583] = 32'b11000001101110000000000000000000;
	assign	vad_gru_input_weights_array[  584] = 32'b11000010110111100000000000000000;
	assign	vad_gru_input_weights_array[  585] = 32'b11000010001010000000000000000000;
	assign	vad_gru_input_weights_array[  586] = 32'b11000010101110100000000000000000;
	assign	vad_gru_input_weights_array[  587] = 32'b11000010111100000000000000000000;
	assign	vad_gru_input_weights_array[  588] = 32'b01000010101101000000000000000000;
	assign	vad_gru_input_weights_array[  589] = 32'b11000010101010100000000000000000;
	assign	vad_gru_input_weights_array[  590] = 32'b11000010010110000000000000000000;
	assign	vad_gru_input_weights_array[  591] = 32'b11000010111011000000000000000000;
	assign	vad_gru_input_weights_array[  592] = 32'b01000010100110000000000000000000;
	assign	vad_gru_input_weights_array[  593] = 32'b11000010100111100000000000000000;
	assign	vad_gru_input_weights_array[  594] = 32'b01000010111110000000000000000000;
	assign	vad_gru_input_weights_array[  595] = 32'b01000010110010100000000000000000;
	assign	vad_gru_input_weights_array[  596] = 32'b11000010100110100000000000000000;
	assign	vad_gru_input_weights_array[  597] = 32'b11000010100101100000000000000000;
	assign	vad_gru_input_weights_array[  598] = 32'b11000001100010000000000000000000;
	assign	vad_gru_input_weights_array[  599] = 32'b11000010100011100000000000000000;
	assign	vad_gru_input_weights_array[  600] = 32'b11000010111001000000000000000000;
	assign	vad_gru_input_weights_array[  601] = 32'b01000010100010000000000000000000;
	assign	vad_gru_input_weights_array[  602] = 32'b01000010010111000000000000000000;
	assign	vad_gru_input_weights_array[  603] = 32'b01000010100111100000000000000000;
	assign	vad_gru_input_weights_array[  604] = 32'b10111111100000000000000000000000;
	assign	vad_gru_input_weights_array[  605] = 32'b11000010111101100000000000000000;
	assign	vad_gru_input_weights_array[  606] = 32'b11000001101000000000000000000000;
	assign	vad_gru_input_weights_array[  607] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  608] = 32'b11000010100000100000000000000000;
	assign	vad_gru_input_weights_array[  609] = 32'b11000010111101100000000000000000;
	assign	vad_gru_input_weights_array[  610] = 32'b11000011000000000000000000000000;
	assign	vad_gru_input_weights_array[  611] = 32'b11000010101011100000000000000000;
	assign	vad_gru_input_weights_array[  612] = 32'b01000010111101100000000000000000;
	assign	vad_gru_input_weights_array[  613] = 32'b01000001000100000000000000000000;
	assign	vad_gru_input_weights_array[  614] = 32'b11000010111001100000000000000000;
	assign	vad_gru_input_weights_array[  615] = 32'b11000001011000000000000000000000;
	assign	vad_gru_input_weights_array[  616] = 32'b01000000111000000000000000000000;
	assign	vad_gru_input_weights_array[  617] = 32'b11000000100000000000000000000000;
	assign	vad_gru_input_weights_array[  618] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  619] = 32'b11000010100111100000000000000000;
	assign	vad_gru_input_weights_array[  620] = 32'b11000010111001100000000000000000;
	assign	vad_gru_input_weights_array[  621] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[  622] = 32'b11000001111000000000000000000000;
	assign	vad_gru_input_weights_array[  623] = 32'b01000010101100100000000000000000;
	assign	vad_gru_input_weights_array[  624] = 32'b11000010101001100000000000000000;
	assign	vad_gru_input_weights_array[  625] = 32'b01000010010001000000000000000000;
	assign	vad_gru_input_weights_array[  626] = 32'b01000010101100100000000000000000;
	assign	vad_gru_input_weights_array[  627] = 32'b01000010111011100000000000000000;
	assign	vad_gru_input_weights_array[  628] = 32'b11000010100010100000000000000000;
	assign	vad_gru_input_weights_array[  629] = 32'b11000000101000000000000000000000;
	assign	vad_gru_input_weights_array[  630] = 32'b01000001010000000000000000000000;
	assign	vad_gru_input_weights_array[  631] = 32'b11000010010001000000000000000000;
	assign	vad_gru_input_weights_array[  632] = 32'b01000010011100000000000000000000;
	assign	vad_gru_input_weights_array[  633] = 32'b01000010011001000000000000000000;
	assign	vad_gru_input_weights_array[  634] = 32'b11000001110000000000000000000000;
	assign	vad_gru_input_weights_array[  635] = 32'b11000010110001100000000000000000;
	assign	vad_gru_input_weights_array[  636] = 32'b11000010110111000000000000000000;
	assign	vad_gru_input_weights_array[  637] = 32'b01000010100110000000000000000000;
	assign	vad_gru_input_weights_array[  638] = 32'b11000010101001100000000000000000;
	assign	vad_gru_input_weights_array[  639] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[  640] = 32'b01000010100100100000000000000000;
	assign	vad_gru_input_weights_array[  641] = 32'b01000010101000100000000000000000;
	assign	vad_gru_input_weights_array[  642] = 32'b01000001001100000000000000000000;
	assign	vad_gru_input_weights_array[  643] = 32'b01000001000000000000000000000000;
	assign	vad_gru_input_weights_array[  644] = 32'b11000010001101000000000000000000;
	assign	vad_gru_input_weights_array[  645] = 32'b00111111100000000000000000000000;
	assign	vad_gru_input_weights_array[  646] = 32'b01000010101001100000000000000000;
	assign	vad_gru_input_weights_array[  647] = 32'b01000001010100000000000000000000;
	assign	vad_gru_input_weights_array[  648] = 32'b11000010100011000000000000000000;
	assign	vad_gru_input_weights_array[  649] = 32'b11000000000000000000000000000000;
	assign	vad_gru_input_weights_array[  650] = 32'b01000010110000100000000000000000;
	assign	vad_gru_input_weights_array[  651] = 32'b01000010111000000000000000000000;
	assign	vad_gru_input_weights_array[  652] = 32'b11000010110000100000000000000000;
	assign	vad_gru_input_weights_array[  653] = 32'b01000010010101000000000000000000;
	assign	vad_gru_input_weights_array[  654] = 32'b11000001000100000000000000000000;
	assign	vad_gru_input_weights_array[  655] = 32'b11000010101111000000000000000000;
	assign	vad_gru_input_weights_array[  656] = 32'b01000010111110000000000000000000;
	assign	vad_gru_input_weights_array[  657] = 32'b01000010001100000000000000000000;
	assign	vad_gru_input_weights_array[  658] = 32'b11000010010001000000000000000000;
	assign	vad_gru_input_weights_array[  659] = 32'b11000001110000000000000000000000;
	assign	vad_gru_input_weights_array[  660] = 32'b01000010010100000000000000000000;
	assign	vad_gru_input_weights_array[  661] = 32'b01000010100110000000000000000000;
	assign	vad_gru_input_weights_array[  662] = 32'b11000010110111000000000000000000;
	assign	vad_gru_input_weights_array[  663] = 32'b11000010100011000000000000000000;
	assign	vad_gru_input_weights_array[  664] = 32'b11000010111001000000000000000000;
	assign	vad_gru_input_weights_array[  665] = 32'b11000001010000000000000000000000;
	assign	vad_gru_input_weights_array[  666] = 32'b01000010100100000000000000000000;
	assign	vad_gru_input_weights_array[  667] = 32'b11000000100000000000000000000000;
	assign	vad_gru_input_weights_array[  668] = 32'b11000010111001000000000000000000;
	assign	vad_gru_input_weights_array[  669] = 32'b01000010001011000000000000000000;
	assign	vad_gru_input_weights_array[  670] = 32'b11000010001011000000000000000000;
	assign	vad_gru_input_weights_array[  671] = 32'b01000010101000100000000000000000;
	assign	vad_gru_input_weights_array[  672] = 32'b01000010110011000000000000000000;
	assign	vad_gru_input_weights_array[  673] = 32'b11000010101010000000000000000000;
	assign	vad_gru_input_weights_array[  674] = 32'b11000001110110000000000000000000;
	assign	vad_gru_input_weights_array[  675] = 32'b01000010011110000000000000000000;
	assign	vad_gru_input_weights_array[  676] = 32'b11000010001000000000000000000000;
	assign	vad_gru_input_weights_array[  677] = 32'b01000010010100000000000000000000;
	assign	vad_gru_input_weights_array[  678] = 32'b01000010011010000000000000000000;
	assign	vad_gru_input_weights_array[  679] = 32'b01000010111110000000000000000000;
	assign	vad_gru_input_weights_array[  680] = 32'b11000010000011000000000000000000;
	assign	vad_gru_input_weights_array[  681] = 32'b11000010010011000000000000000000;
	assign	vad_gru_input_weights_array[  682] = 32'b11000010111101100000000000000000;
	assign	vad_gru_input_weights_array[  683] = 32'b11000010001011000000000000000000;
	assign	vad_gru_input_weights_array[  684] = 32'b01000010011000000000000000000000;
	assign	vad_gru_input_weights_array[  685] = 32'b11000010100101100000000000000000;
	assign	vad_gru_input_weights_array[  686] = 32'b11000010000010000000000000000000;
	assign	vad_gru_input_weights_array[  687] = 32'b11000010000011000000000000000000;
	assign	vad_gru_input_weights_array[  688] = 32'b11000010110101000000000000000000;
	assign	vad_gru_input_weights_array[  689] = 32'b01000010101110100000000000000000;
	assign	vad_gru_input_weights_array[  690] = 32'b11000010001011000000000000000000;
	assign	vad_gru_input_weights_array[  691] = 32'b01000001011000000000000000000000;
	assign	vad_gru_input_weights_array[  692] = 32'b11000001100000000000000000000000;
	assign	vad_gru_input_weights_array[  693] = 32'b01000010001110000000000000000000;
	assign	vad_gru_input_weights_array[  694] = 32'b01000010011110000000000000000000;
	assign	vad_gru_input_weights_array[  695] = 32'b11000010110000100000000000000000;
	assign	vad_gru_input_weights_array[  696] = 32'b01000001101010000000000000000000;
	assign	vad_gru_input_weights_array[  697] = 32'b01000001111100000000000000000000;
	assign	vad_gru_input_weights_array[  698] = 32'b11000010010101000000000000000000;
	assign	vad_gru_input_weights_array[  699] = 32'b01000001101010000000000000000000;
	assign	vad_gru_input_weights_array[  700] = 32'b11000001001100000000000000000000;
	assign	vad_gru_input_weights_array[  701] = 32'b11000010000001000000000000000000;
	assign	vad_gru_input_weights_array[  702] = 32'b11000001101000000000000000000000;
	assign	vad_gru_input_weights_array[  703] = 32'b11000010101111100000000000000000;
	assign	vad_gru_input_weights_array[  704] = 32'b01000000100000000000000000000000;
	assign	vad_gru_input_weights_array[  705] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  706] = 32'b01000001010000000000000000000000;
	assign	vad_gru_input_weights_array[  707] = 32'b01000010001101000000000000000000;
	assign	vad_gru_input_weights_array[  708] = 32'b01000001101000000000000000000000;
	assign	vad_gru_input_weights_array[  709] = 32'b01000010110110000000000000000000;
	assign	vad_gru_input_weights_array[  710] = 32'b01000010101010100000000000000000;
	assign	vad_gru_input_weights_array[  711] = 32'b01000001001100000000000000000000;
	assign	vad_gru_input_weights_array[  712] = 32'b01000001101000000000000000000000;
	assign	vad_gru_input_weights_array[  713] = 32'b11000010001000000000000000000000;
	assign	vad_gru_input_weights_array[  714] = 32'b01000010110001100000000000000000;
	assign	vad_gru_input_weights_array[  715] = 32'b01000000100000000000000000000000;
	assign	vad_gru_input_weights_array[  716] = 32'b11000001110010000000000000000000;
	assign	vad_gru_input_weights_array[  717] = 32'b11000001100100000000000000000000;
	assign	vad_gru_input_weights_array[  718] = 32'b11000001101110000000000000000000;
	assign	vad_gru_input_weights_array[  719] = 32'b11000001010000000000000000000000;
	assign	vad_gru_input_weights_array[  720] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  721] = 32'b11000010010111000000000000000000;
	assign	vad_gru_input_weights_array[  722] = 32'b11000001101000000000000000000000;
	assign	vad_gru_input_weights_array[  723] = 32'b11000010001100000000000000000000;
	assign	vad_gru_input_weights_array[  724] = 32'b11000010010011000000000000000000;
	assign	vad_gru_input_weights_array[  725] = 32'b01000010101101100000000000000000;
	assign	vad_gru_input_weights_array[  726] = 32'b11000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  727] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  728] = 32'b11000010001100000000000000000000;
	assign	vad_gru_input_weights_array[  729] = 32'b01000000111000000000000000000000;
	assign	vad_gru_input_weights_array[  730] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  731] = 32'b01000010100111000000000000000000;
	assign	vad_gru_input_weights_array[  732] = 32'b01000010000110000000000000000000;
	assign	vad_gru_input_weights_array[  733] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[  734] = 32'b11000000110000000000000000000000;
	assign	vad_gru_input_weights_array[  735] = 32'b11000010101111000000000000000000;
	assign	vad_gru_input_weights_array[  736] = 32'b11000010110011100000000000000000;
	assign	vad_gru_input_weights_array[  737] = 32'b01000010100100100000000000000000;
	assign	vad_gru_input_weights_array[  738] = 32'b01000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  739] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  740] = 32'b01000001100100000000000000000000;
	assign	vad_gru_input_weights_array[  741] = 32'b01000010011011000000000000000000;
	assign	vad_gru_input_weights_array[  742] = 32'b11000010001110000000000000000000;
	assign	vad_gru_input_weights_array[  743] = 32'b01000010110101000000000000000000;
	assign	vad_gru_input_weights_array[  744] = 32'b01000010100110000000000000000000;
	assign	vad_gru_input_weights_array[  745] = 32'b01000010111010000000000000000000;
	assign	vad_gru_input_weights_array[  746] = 32'b11000001111110000000000000000000;
	assign	vad_gru_input_weights_array[  747] = 32'b01000010100101100000000000000000;
	assign	vad_gru_input_weights_array[  748] = 32'b11000000100000000000000000000000;
	assign	vad_gru_input_weights_array[  749] = 32'b01000010101110000000000000000000;
	assign	vad_gru_input_weights_array[  750] = 32'b01000010110011000000000000000000;
	assign	vad_gru_input_weights_array[  751] = 32'b01000010000000000000000000000000;
	assign	vad_gru_input_weights_array[  752] = 32'b11000001111110000000000000000000;
	assign	vad_gru_input_weights_array[  753] = 32'b01000010100100100000000000000000;
	assign	vad_gru_input_weights_array[  754] = 32'b01000010001010000000000000000000;
	assign	vad_gru_input_weights_array[  755] = 32'b11000001101010000000000000000000;
	assign	vad_gru_input_weights_array[  756] = 32'b11000001111000000000000000000000;
	assign	vad_gru_input_weights_array[  757] = 32'b01000010011001000000000000000000;
	assign	vad_gru_input_weights_array[  758] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  759] = 32'b11000001000000000000000000000000;
	assign	vad_gru_input_weights_array[  760] = 32'b11000010110101100000000000000000;
	assign	vad_gru_input_weights_array[  761] = 32'b01000010111001100000000000000000;
	assign	vad_gru_input_weights_array[  762] = 32'b01000010111110000000000000000000;
	assign	vad_gru_input_weights_array[  763] = 32'b11000010101111000000000000000000;
	assign	vad_gru_input_weights_array[  764] = 32'b11000000100000000000000000000000;
	assign	vad_gru_input_weights_array[  765] = 32'b11000011000000000000000000000000;
	assign	vad_gru_input_weights_array[  766] = 32'b01000001111010000000000000000000;
	assign	vad_gru_input_weights_array[  767] = 32'b11000010011001000000000000000000;
	assign	vad_gru_input_weights_array[  768] = 32'b01000010100011000000000000000000;
	assign	vad_gru_input_weights_array[  769] = 32'b11000010101001000000000000000000;
	assign	vad_gru_input_weights_array[  770] = 32'b01000010010010000000000000000000;
	assign	vad_gru_input_weights_array[  771] = 32'b11000001010100000000000000000000;
	assign	vad_gru_input_weights_array[  772] = 32'b11000010001100000000000000000000;
	assign	vad_gru_input_weights_array[  773] = 32'b01000010000110000000000000000000;
	assign	vad_gru_input_weights_array[  774] = 32'b01000010100001100000000000000000;
	assign	vad_gru_input_weights_array[  775] = 32'b11000010101110100000000000000000;
	assign	vad_gru_input_weights_array[  776] = 32'b01000000110000000000000000000000;
	assign	vad_gru_input_weights_array[  777] = 32'b11000010000111000000000000000000;
	assign	vad_gru_input_weights_array[  778] = 32'b11000010001110000000000000000000;
	assign	vad_gru_input_weights_array[  779] = 32'b01000010011000000000000000000000;
	assign	vad_gru_input_weights_array[  780] = 32'b01000010100010000000000000000000;
	assign	vad_gru_input_weights_array[  781] = 32'b01000001110110000000000000000000;
	assign	vad_gru_input_weights_array[  782] = 32'b01000010011101000000000000000000;
	assign	vad_gru_input_weights_array[  783] = 32'b01000001110100000000000000000000;
	assign	vad_gru_input_weights_array[  784] = 32'b01000001100100000000000000000000;
	assign	vad_gru_input_weights_array[  785] = 32'b11000010100100000000000000000000;
	assign	vad_gru_input_weights_array[  786] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  787] = 32'b01000001101100000000000000000000;
	assign	vad_gru_input_weights_array[  788] = 32'b01000001100100000000000000000000;
	assign	vad_gru_input_weights_array[  789] = 32'b11000001111110000000000000000000;
	assign	vad_gru_input_weights_array[  790] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  791] = 32'b01000010011101000000000000000000;
	assign	vad_gru_input_weights_array[  792] = 32'b11000010100000100000000000000000;
	assign	vad_gru_input_weights_array[  793] = 32'b11000010000110000000000000000000;
	assign	vad_gru_input_weights_array[  794] = 32'b00111111100000000000000000000000;
	assign	vad_gru_input_weights_array[  795] = 32'b11000010100001100000000000000000;
	assign	vad_gru_input_weights_array[  796] = 32'b10111111100000000000000000000000;
	assign	vad_gru_input_weights_array[  797] = 32'b01000001000000000000000000000000;
	assign	vad_gru_input_weights_array[  798] = 32'b11000010100100100000000000000000;
	assign	vad_gru_input_weights_array[  799] = 32'b01000010001110000000000000000000;
	assign	vad_gru_input_weights_array[  800] = 32'b11000010111010000000000000000000;
	assign	vad_gru_input_weights_array[  801] = 32'b11000010101111000000000000000000;
	assign	vad_gru_input_weights_array[  802] = 32'b01000010011010000000000000000000;
	assign	vad_gru_input_weights_array[  803] = 32'b11000010010001000000000000000000;
	assign	vad_gru_input_weights_array[  804] = 32'b01000010100011100000000000000000;
	assign	vad_gru_input_weights_array[  805] = 32'b11000010001000000000000000000000;
	assign	vad_gru_input_weights_array[  806] = 32'b11000010011111000000000000000000;
	assign	vad_gru_input_weights_array[  807] = 32'b11000010101001000000000000000000;
	assign	vad_gru_input_weights_array[  808] = 32'b11000001101000000000000000000000;
	assign	vad_gru_input_weights_array[  809] = 32'b11000010011100000000000000000000;
	assign	vad_gru_input_weights_array[  810] = 32'b01000010101110100000000000000000;
	assign	vad_gru_input_weights_array[  811] = 32'b01000010100110000000000000000000;
	assign	vad_gru_input_weights_array[  812] = 32'b01000010100010100000000000000000;
	assign	vad_gru_input_weights_array[  813] = 32'b11000010110101000000000000000000;
	assign	vad_gru_input_weights_array[  814] = 32'b01000010000010000000000000000000;
	assign	vad_gru_input_weights_array[  815] = 32'b11000001111110000000000000000000;
	assign	vad_gru_input_weights_array[  816] = 32'b01000000100000000000000000000000;
	assign	vad_gru_input_weights_array[  817] = 32'b11000001110010000000000000000000;
	assign	vad_gru_input_weights_array[  818] = 32'b01000010110101100000000000000000;
	assign	vad_gru_input_weights_array[  819] = 32'b11000001100100000000000000000000;
	assign	vad_gru_input_weights_array[  820] = 32'b01000010001101000000000000000000;
	assign	vad_gru_input_weights_array[  821] = 32'b01000000100000000000000000000000;
	assign	vad_gru_input_weights_array[  822] = 32'b11000010011101000000000000000000;
	assign	vad_gru_input_weights_array[  823] = 32'b01000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  824] = 32'b01000010010110000000000000000000;
	assign	vad_gru_input_weights_array[  825] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  826] = 32'b11000010111110100000000000000000;
	assign	vad_gru_input_weights_array[  827] = 32'b01000010001001000000000000000000;
	assign	vad_gru_input_weights_array[  828] = 32'b01000001100110000000000000000000;
	assign	vad_gru_input_weights_array[  829] = 32'b01000010001100000000000000000000;
	assign	vad_gru_input_weights_array[  830] = 32'b01000010000000000000000000000000;
	assign	vad_gru_input_weights_array[  831] = 32'b11000010110001000000000000000000;
	assign	vad_gru_input_weights_array[  832] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[  833] = 32'b11000001110000000000000000000000;
	assign	vad_gru_input_weights_array[  834] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[  835] = 32'b11000010110000000000000000000000;
	assign	vad_gru_input_weights_array[  836] = 32'b11000010111110100000000000000000;
	assign	vad_gru_input_weights_array[  837] = 32'b01000001011100000000000000000000;
	assign	vad_gru_input_weights_array[  838] = 32'b01000010101011100000000000000000;
	assign	vad_gru_input_weights_array[  839] = 32'b11000000100000000000000000000000;
	assign	vad_gru_input_weights_array[  840] = 32'b11000010101101000000000000000000;
	assign	vad_gru_input_weights_array[  841] = 32'b01000001100100000000000000000000;
	assign	vad_gru_input_weights_array[  842] = 32'b11000010001000000000000000000000;
	assign	vad_gru_input_weights_array[  843] = 32'b01000001111000000000000000000000;
	assign	vad_gru_input_weights_array[  844] = 32'b11000010100010100000000000000000;
	assign	vad_gru_input_weights_array[  845] = 32'b01000010100001100000000000000000;
	assign	vad_gru_input_weights_array[  846] = 32'b01000001101100000000000000000000;
	assign	vad_gru_input_weights_array[  847] = 32'b01000010001001000000000000000000;
	assign	vad_gru_input_weights_array[  848] = 32'b01000010000111000000000000000000;
	assign	vad_gru_input_weights_array[  849] = 32'b01000000111000000000000000000000;
	assign	vad_gru_input_weights_array[  850] = 32'b11000010010000000000000000000000;
	assign	vad_gru_input_weights_array[  851] = 32'b11000010001100000000000000000000;
	assign	vad_gru_input_weights_array[  852] = 32'b01000001010000000000000000000000;
	assign	vad_gru_input_weights_array[  853] = 32'b01000010100010100000000000000000;
	assign	vad_gru_input_weights_array[  854] = 32'b11000001010100000000000000000000;
	assign	vad_gru_input_weights_array[  855] = 32'b01000000000000000000000000000000;
	assign	vad_gru_input_weights_array[  856] = 32'b01000010001100000000000000000000;
	assign	vad_gru_input_weights_array[  857] = 32'b11000010000110000000000000000000;
	assign	vad_gru_input_weights_array[  858] = 32'b01000010110111100000000000000000;
	assign	vad_gru_input_weights_array[  859] = 32'b11000000111000000000000000000000;
	assign	vad_gru_input_weights_array[  860] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  861] = 32'b11000001101100000000000000000000;
	assign	vad_gru_input_weights_array[  862] = 32'b11000001000100000000000000000000;
	assign	vad_gru_input_weights_array[  863] = 32'b01000010100101000000000000000000;
	assign	vad_gru_input_weights_array[  864] = 32'b11000011000000000000000000000000;
	assign	vad_gru_input_weights_array[  865] = 32'b11000010000100000000000000000000;
	assign	vad_gru_input_weights_array[  866] = 32'b11000000111000000000000000000000;
	assign	vad_gru_input_weights_array[  867] = 32'b11000010111101100000000000000000;
	assign	vad_gru_input_weights_array[  868] = 32'b11000001011100000000000000000000;
	assign	vad_gru_input_weights_array[  869] = 32'b11000010100111100000000000000000;
	assign	vad_gru_input_weights_array[  870] = 32'b11000010101101100000000000000000;
	assign	vad_gru_input_weights_array[  871] = 32'b11000010000101000000000000000000;
	assign	vad_gru_input_weights_array[  872] = 32'b11000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  873] = 32'b11000010111101000000000000000000;
	assign	vad_gru_input_weights_array[  874] = 32'b01000010110100000000000000000000;
	assign	vad_gru_input_weights_array[  875] = 32'b01000001111100000000000000000000;
	assign	vad_gru_input_weights_array[  876] = 32'b01000000111000000000000000000000;
	assign	vad_gru_input_weights_array[  877] = 32'b01000010110001000000000000000000;
	assign	vad_gru_input_weights_array[  878] = 32'b11000010000101000000000000000000;
	assign	vad_gru_input_weights_array[  879] = 32'b01000010110111100000000000000000;
	assign	vad_gru_input_weights_array[  880] = 32'b11000010111010000000000000000000;
	assign	vad_gru_input_weights_array[  881] = 32'b11000010001111000000000000000000;
	assign	vad_gru_input_weights_array[  882] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  883] = 32'b11000010001101000000000000000000;
	assign	vad_gru_input_weights_array[  884] = 32'b01000010111011000000000000000000;
	assign	vad_gru_input_weights_array[  885] = 32'b11000010110111100000000000000000;
	assign	vad_gru_input_weights_array[  886] = 32'b11000010111101100000000000000000;
	assign	vad_gru_input_weights_array[  887] = 32'b11000010111100000000000000000000;
	assign	vad_gru_input_weights_array[  888] = 32'b11000010100110100000000000000000;
	assign	vad_gru_input_weights_array[  889] = 32'b11000010100000000000000000000000;
	assign	vad_gru_input_weights_array[  890] = 32'b11000010111110100000000000000000;
	assign	vad_gru_input_weights_array[  891] = 32'b01000010111110000000000000000000;
	assign	vad_gru_input_weights_array[  892] = 32'b01000010100110100000000000000000;
	assign	vad_gru_input_weights_array[  893] = 32'b01000010110111100000000000000000;
	assign	vad_gru_input_weights_array[  894] = 32'b01000010100110100000000000000000;
	assign	vad_gru_input_weights_array[  895] = 32'b01000001100100000000000000000000;
	assign	vad_gru_input_weights_array[  896] = 32'b11000010111000100000000000000000;
	assign	vad_gru_input_weights_array[  897] = 32'b01000010111010100000000000000000;
	assign	vad_gru_input_weights_array[  898] = 32'b11000001000100000000000000000000;
	assign	vad_gru_input_weights_array[  899] = 32'b01000010100001100000000000000000;
	assign	vad_gru_input_weights_array[  900] = 32'b11000010100110100000000000000000;
	assign	vad_gru_input_weights_array[  901] = 32'b01000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  902] = 32'b01000010010001000000000000000000;
	assign	vad_gru_input_weights_array[  903] = 32'b11000001101000000000000000000000;
	assign	vad_gru_input_weights_array[  904] = 32'b11000010111110000000000000000000;
	assign	vad_gru_input_weights_array[  905] = 32'b01000010000111000000000000000000;
	assign	vad_gru_input_weights_array[  906] = 32'b01000010001001000000000000000000;
	assign	vad_gru_input_weights_array[  907] = 32'b11000010111110000000000000000000;
	assign	vad_gru_input_weights_array[  908] = 32'b11000010000010000000000000000000;
	assign	vad_gru_input_weights_array[  909] = 32'b01000010111001000000000000000000;
	assign	vad_gru_input_weights_array[  910] = 32'b11000010101011100000000000000000;
	assign	vad_gru_input_weights_array[  911] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  912] = 32'b01000010110001000000000000000000;
	assign	vad_gru_input_weights_array[  913] = 32'b11000001101000000000000000000000;
	assign	vad_gru_input_weights_array[  914] = 32'b01000010011011000000000000000000;
	assign	vad_gru_input_weights_array[  915] = 32'b11000001100010000000000000000000;
	assign	vad_gru_input_weights_array[  916] = 32'b11000001110000000000000000000000;
	assign	vad_gru_input_weights_array[  917] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[  918] = 32'b01000010110101100000000000000000;
	assign	vad_gru_input_weights_array[  919] = 32'b01000010010110000000000000000000;
	assign	vad_gru_input_weights_array[  920] = 32'b01000010000011000000000000000000;
	assign	vad_gru_input_weights_array[  921] = 32'b01000010000001000000000000000000;
	assign	vad_gru_input_weights_array[  922] = 32'b11000010001100000000000000000000;
	assign	vad_gru_input_weights_array[  923] = 32'b01000001010000000000000000000000;
	assign	vad_gru_input_weights_array[  924] = 32'b11000001111010000000000000000000;
	assign	vad_gru_input_weights_array[  925] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[  926] = 32'b11000010100011100000000000000000;
	assign	vad_gru_input_weights_array[  927] = 32'b11000001111000000000000000000000;
	assign	vad_gru_input_weights_array[  928] = 32'b11000010011111000000000000000000;
	assign	vad_gru_input_weights_array[  929] = 32'b11000010111001000000000000000000;
	assign	vad_gru_input_weights_array[  930] = 32'b01000001111000000000000000000000;
	assign	vad_gru_input_weights_array[  931] = 32'b11000001100010000000000000000000;
	assign	vad_gru_input_weights_array[  932] = 32'b01000010111100100000000000000000;
	assign	vad_gru_input_weights_array[  933] = 32'b11000010000100000000000000000000;
	assign	vad_gru_input_weights_array[  934] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  935] = 32'b01000010101100100000000000000000;
	assign	vad_gru_input_weights_array[  936] = 32'b11000010111101000000000000000000;
	assign	vad_gru_input_weights_array[  937] = 32'b11000010010001000000000000000000;
	assign	vad_gru_input_weights_array[  938] = 32'b11000001100100000000000000000000;
	assign	vad_gru_input_weights_array[  939] = 32'b11000010010000000000000000000000;
	assign	vad_gru_input_weights_array[  940] = 32'b01000001100010000000000000000000;
	assign	vad_gru_input_weights_array[  941] = 32'b01000001110000000000000000000000;
	assign	vad_gru_input_weights_array[  942] = 32'b01000001100110000000000000000000;
	assign	vad_gru_input_weights_array[  943] = 32'b11000010100000000000000000000000;
	assign	vad_gru_input_weights_array[  944] = 32'b11000011000000000000000000000000;
	assign	vad_gru_input_weights_array[  945] = 32'b01000001010100000000000000000000;
	assign	vad_gru_input_weights_array[  946] = 32'b01000010101011000000000000000000;
	assign	vad_gru_input_weights_array[  947] = 32'b01000010001101000000000000000000;
	assign	vad_gru_input_weights_array[  948] = 32'b01000001010100000000000000000000;
	assign	vad_gru_input_weights_array[  949] = 32'b11000010010001000000000000000000;
	assign	vad_gru_input_weights_array[  950] = 32'b01000010010111000000000000000000;
	assign	vad_gru_input_weights_array[  951] = 32'b01000010101010000000000000000000;
	assign	vad_gru_input_weights_array[  952] = 32'b01000010010000000000000000000000;
	assign	vad_gru_input_weights_array[  953] = 32'b01000010101000000000000000000000;
	assign	vad_gru_input_weights_array[  954] = 32'b11000010000111000000000000000000;
	assign	vad_gru_input_weights_array[  955] = 32'b01000010110001100000000000000000;
	assign	vad_gru_input_weights_array[  956] = 32'b11000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  957] = 32'b01000010100011000000000000000000;
	assign	vad_gru_input_weights_array[  958] = 32'b11000010000001000000000000000000;
	assign	vad_gru_input_weights_array[  959] = 32'b01000001111100000000000000000000;
	assign	vad_gru_input_weights_array[  960] = 32'b01000010010010000000000000000000;
	assign	vad_gru_input_weights_array[  961] = 32'b01000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  962] = 32'b11000010100000100000000000000000;
	assign	vad_gru_input_weights_array[  963] = 32'b11000010111010100000000000000000;
	assign	vad_gru_input_weights_array[  964] = 32'b11000001010100000000000000000000;
	assign	vad_gru_input_weights_array[  965] = 32'b11000001101000000000000000000000;
	assign	vad_gru_input_weights_array[  966] = 32'b11000001110000000000000000000000;
	assign	vad_gru_input_weights_array[  967] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[  968] = 32'b01000010111001100000000000000000;
	assign	vad_gru_input_weights_array[  969] = 32'b11000010100100000000000000000000;
	assign	vad_gru_input_weights_array[  970] = 32'b11000010110100000000000000000000;
	assign	vad_gru_input_weights_array[  971] = 32'b01000010011111000000000000000000;
	assign	vad_gru_input_weights_array[  972] = 32'b01000010111111000000000000000000;
	assign	vad_gru_input_weights_array[  973] = 32'b11000010001010000000000000000000;
	assign	vad_gru_input_weights_array[  974] = 32'b01000010011001000000000000000000;
	assign	vad_gru_input_weights_array[  975] = 32'b01000001100010000000000000000000;
	assign	vad_gru_input_weights_array[  976] = 32'b01000010001110000000000000000000;
	assign	vad_gru_input_weights_array[  977] = 32'b01000001101010000000000000000000;
	assign	vad_gru_input_weights_array[  978] = 32'b01000010111011100000000000000000;
	assign	vad_gru_input_weights_array[  979] = 32'b01000010110111000000000000000000;
	assign	vad_gru_input_weights_array[  980] = 32'b11000010110010000000000000000000;
	assign	vad_gru_input_weights_array[  981] = 32'b11000010011100000000000000000000;
	assign	vad_gru_input_weights_array[  982] = 32'b11000010111000000000000000000000;
	assign	vad_gru_input_weights_array[  983] = 32'b01000010011110000000000000000000;
	assign	vad_gru_input_weights_array[  984] = 32'b11000010000001000000000000000000;
	assign	vad_gru_input_weights_array[  985] = 32'b01000001111000000000000000000000;
	assign	vad_gru_input_weights_array[  986] = 32'b01000001110100000000000000000000;
	assign	vad_gru_input_weights_array[  987] = 32'b11000001101100000000000000000000;
	assign	vad_gru_input_weights_array[  988] = 32'b11000010011100000000000000000000;
	assign	vad_gru_input_weights_array[  989] = 32'b11000010000001000000000000000000;
	assign	vad_gru_input_weights_array[  990] = 32'b11000010010110000000000000000000;
	assign	vad_gru_input_weights_array[  991] = 32'b01000010100111000000000000000000;
	assign	vad_gru_input_weights_array[  992] = 32'b01000001110010000000000000000000;
	assign	vad_gru_input_weights_array[  993] = 32'b01000010000000000000000000000000;
	assign	vad_gru_input_weights_array[  994] = 32'b11000010111001000000000000000000;
	assign	vad_gru_input_weights_array[  995] = 32'b01000010101011000000000000000000;
	assign	vad_gru_input_weights_array[  996] = 32'b01000010001100000000000000000000;
	assign	vad_gru_input_weights_array[  997] = 32'b01000001110100000000000000000000;
	assign	vad_gru_input_weights_array[  998] = 32'b01000010001011000000000000000000;
	assign	vad_gru_input_weights_array[  999] = 32'b01000010100110000000000000000000;
	assign	vad_gru_input_weights_array[ 1000] = 32'b01000010111100100000000000000000;
	assign	vad_gru_input_weights_array[ 1001] = 32'b01000001100110000000000000000000;
	assign	vad_gru_input_weights_array[ 1002] = 32'b01000010110000100000000000000000;
	assign	vad_gru_input_weights_array[ 1003] = 32'b11000000000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1004] = 32'b11000000010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1005] = 32'b11000010100100100000000000000000;
	assign	vad_gru_input_weights_array[ 1006] = 32'b11000010100010000000000000000000;
	assign	vad_gru_input_weights_array[ 1007] = 32'b01000000110000000000000000000000;
	assign	vad_gru_input_weights_array[ 1008] = 32'b11000010111010000000000000000000;
	assign	vad_gru_input_weights_array[ 1009] = 32'b01000000110000000000000000000000;
	assign	vad_gru_input_weights_array[ 1010] = 32'b11000010001011000000000000000000;
	assign	vad_gru_input_weights_array[ 1011] = 32'b11000010110000100000000000000000;
	assign	vad_gru_input_weights_array[ 1012] = 32'b01000010001110000000000000000000;
	assign	vad_gru_input_weights_array[ 1013] = 32'b11000011000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1014] = 32'b11000010111100000000000000000000;
	assign	vad_gru_input_weights_array[ 1015] = 32'b11000001111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1016] = 32'b11000010111011100000000000000000;
	assign	vad_gru_input_weights_array[ 1017] = 32'b11000001111010000000000000000000;
	assign	vad_gru_input_weights_array[ 1018] = 32'b01000001100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1019] = 32'b01000001100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1020] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[ 1021] = 32'b11000011000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1022] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[ 1023] = 32'b11000010001110000000000000000000;
	assign	vad_gru_input_weights_array[ 1024] = 32'b11000001000100000000000000000000;
	assign	vad_gru_input_weights_array[ 1025] = 32'b11000000010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1026] = 32'b01000010101110000000000000000000;
	assign	vad_gru_input_weights_array[ 1027] = 32'b11000001111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1028] = 32'b11000010100110000000000000000000;
	assign	vad_gru_input_weights_array[ 1029] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[ 1030] = 32'b11000000010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1031] = 32'b11000010110101100000000000000000;
	assign	vad_gru_input_weights_array[ 1032] = 32'b11000001010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1033] = 32'b11000001101110000000000000000000;
	assign	vad_gru_input_weights_array[ 1034] = 32'b11000010100010100000000000000000;
	assign	vad_gru_input_weights_array[ 1035] = 32'b01000000101000000000000000000000;
	assign	vad_gru_input_weights_array[ 1036] = 32'b01000010010011000000000000000000;
	assign	vad_gru_input_weights_array[ 1037] = 32'b01000001110110000000000000000000;
	assign	vad_gru_input_weights_array[ 1038] = 32'b11000010001010000000000000000000;
	assign	vad_gru_input_weights_array[ 1039] = 32'b01000001101110000000000000000000;
	assign	vad_gru_input_weights_array[ 1040] = 32'b11000010100011000000000000000000;
	assign	vad_gru_input_weights_array[ 1041] = 32'b11000011000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1042] = 32'b11000001111010000000000000000000;
	assign	vad_gru_input_weights_array[ 1043] = 32'b01000001101100000000000000000000;
	assign	vad_gru_input_weights_array[ 1044] = 32'b01000001111010000000000000000000;
	assign	vad_gru_input_weights_array[ 1045] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[ 1046] = 32'b11000010010111000000000000000000;
	assign	vad_gru_input_weights_array[ 1047] = 32'b01000010010010000000000000000000;
	assign	vad_gru_input_weights_array[ 1048] = 32'b11000010100011100000000000000000;
	assign	vad_gru_input_weights_array[ 1049] = 32'b11000000010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1050] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[ 1051] = 32'b01000010001100000000000000000000;
	assign	vad_gru_input_weights_array[ 1052] = 32'b11000001110110000000000000000000;
	assign	vad_gru_input_weights_array[ 1053] = 32'b11000010100011000000000000000000;
	assign	vad_gru_input_weights_array[ 1054] = 32'b11000010011111000000000000000000;
	assign	vad_gru_input_weights_array[ 1055] = 32'b11000010100001000000000000000000;
	assign	vad_gru_input_weights_array[ 1056] = 32'b11000010100011000000000000000000;
	assign	vad_gru_input_weights_array[ 1057] = 32'b01000010110100000000000000000000;
	assign	vad_gru_input_weights_array[ 1058] = 32'b01000010101011000000000000000000;
	assign	vad_gru_input_weights_array[ 1059] = 32'b01000010111001100000000000000000;
	assign	vad_gru_input_weights_array[ 1060] = 32'b01000001111010000000000000000000;
	assign	vad_gru_input_weights_array[ 1061] = 32'b11000010101110000000000000000000;
	assign	vad_gru_input_weights_array[ 1062] = 32'b01000010001001000000000000000000;
	assign	vad_gru_input_weights_array[ 1063] = 32'b11000010101101000000000000000000;
	assign	vad_gru_input_weights_array[ 1064] = 32'b01000010001100000000000000000000;
	assign	vad_gru_input_weights_array[ 1065] = 32'b11000001001100000000000000000000;
	assign	vad_gru_input_weights_array[ 1066] = 32'b11000001111000000000000000000000;
	assign	vad_gru_input_weights_array[ 1067] = 32'b01000001101000000000000000000000;
	assign	vad_gru_input_weights_array[ 1068] = 32'b11000001001100000000000000000000;
	assign	vad_gru_input_weights_array[ 1069] = 32'b11000010011111000000000000000000;
	assign	vad_gru_input_weights_array[ 1070] = 32'b11000001100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1071] = 32'b01000010001011000000000000000000;
	assign	vad_gru_input_weights_array[ 1072] = 32'b01000001111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1073] = 32'b01000001100010000000000000000000;
	assign	vad_gru_input_weights_array[ 1074] = 32'b11000010100100100000000000000000;
	assign	vad_gru_input_weights_array[ 1075] = 32'b11000001111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1076] = 32'b10111111100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1077] = 32'b11000001100010000000000000000000;
	assign	vad_gru_input_weights_array[ 1078] = 32'b11000001001100000000000000000000;
	assign	vad_gru_input_weights_array[ 1079] = 32'b11000010000111000000000000000000;
	assign	vad_gru_input_weights_array[ 1080] = 32'b01000010011000000000000000000000;
	assign	vad_gru_input_weights_array[ 1081] = 32'b01000001100100000000000000000000;
	assign	vad_gru_input_weights_array[ 1082] = 32'b01000010111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1083] = 32'b01000010100100000000000000000000;
	assign	vad_gru_input_weights_array[ 1084] = 32'b11000001011000000000000000000000;
	assign	vad_gru_input_weights_array[ 1085] = 32'b01000001111000000000000000000000;
	assign	vad_gru_input_weights_array[ 1086] = 32'b01000010100010100000000000000000;
	assign	vad_gru_input_weights_array[ 1087] = 32'b11000010111100100000000000000000;
	assign	vad_gru_input_weights_array[ 1088] = 32'b11000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1089] = 32'b01000010000010000000000000000000;
	assign	vad_gru_input_weights_array[ 1090] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[ 1091] = 32'b01000010011111000000000000000000;
	assign	vad_gru_input_weights_array[ 1092] = 32'b01000010101011000000000000000000;
	assign	vad_gru_input_weights_array[ 1093] = 32'b11000010101000000000000000000000;
	assign	vad_gru_input_weights_array[ 1094] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[ 1095] = 32'b11000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1096] = 32'b11000010111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1097] = 32'b11000010001111000000000000000000;
	assign	vad_gru_input_weights_array[ 1098] = 32'b01000010111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1099] = 32'b01000010100110100000000000000000;
	assign	vad_gru_input_weights_array[ 1100] = 32'b01000010111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1101] = 32'b11000001100110000000000000000000;
	assign	vad_gru_input_weights_array[ 1102] = 32'b01000001101110000000000000000000;
	assign	vad_gru_input_weights_array[ 1103] = 32'b11000000111000000000000000000000;
	assign	vad_gru_input_weights_array[ 1104] = 32'b11000010010010000000000000000000;
	assign	vad_gru_input_weights_array[ 1105] = 32'b01000010110000000000000000000000;
	assign	vad_gru_input_weights_array[ 1106] = 32'b11000011000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1107] = 32'b11000010101110100000000000000000;
	assign	vad_gru_input_weights_array[ 1108] = 32'b01000010110011000000000000000000;
	assign	vad_gru_input_weights_array[ 1109] = 32'b11000010010101000000000000000000;
	assign	vad_gru_input_weights_array[ 1110] = 32'b11000010000100000000000000000000;
	assign	vad_gru_input_weights_array[ 1111] = 32'b11000010101011100000000000000000;
	assign	vad_gru_input_weights_array[ 1112] = 32'b01000010111011100000000000000000;
	assign	vad_gru_input_weights_array[ 1113] = 32'b11000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1114] = 32'b01000010101110000000000000000000;
	assign	vad_gru_input_weights_array[ 1115] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[ 1116] = 32'b01000010111011000000000000000000;
	assign	vad_gru_input_weights_array[ 1117] = 32'b01000010110011000000000000000000;
	assign	vad_gru_input_weights_array[ 1118] = 32'b01000010100100000000000000000000;
	assign	vad_gru_input_weights_array[ 1119] = 32'b11000000000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1120] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1121] = 32'b01000001001000000000000000000000;
	assign	vad_gru_input_weights_array[ 1122] = 32'b01000010110000100000000000000000;
	assign	vad_gru_input_weights_array[ 1123] = 32'b01000010111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1124] = 32'b11000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1125] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1126] = 32'b01000010100011100000000000000000;
	assign	vad_gru_input_weights_array[ 1127] = 32'b11000001101000000000000000000000;
	assign	vad_gru_input_weights_array[ 1128] = 32'b11000010001111000000000000000000;
	assign	vad_gru_input_weights_array[ 1129] = 32'b11000010111010000000000000000000;
	assign	vad_gru_input_weights_array[ 1130] = 32'b11000010111100100000000000000000;
	assign	vad_gru_input_weights_array[ 1131] = 32'b11000000100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1132] = 32'b11000001000100000000000000000000;
	assign	vad_gru_input_weights_array[ 1133] = 32'b11000010000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1134] = 32'b01000010100111100000000000000000;
	assign	vad_gru_input_weights_array[ 1135] = 32'b11000010111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1136] = 32'b11000010000100000000000000000000;
	assign	vad_gru_input_weights_array[ 1137] = 32'b01000010000001000000000000000000;
	assign	vad_gru_input_weights_array[ 1138] = 32'b11000011000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1139] = 32'b11000010100101000000000000000000;
	assign	vad_gru_input_weights_array[ 1140] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1141] = 32'b01000001101110000000000000000000;
	assign	vad_gru_input_weights_array[ 1142] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[ 1143] = 32'b11000001111010000000000000000000;
	assign	vad_gru_input_weights_array[ 1144] = 32'b11000010111001100000000000000000;
	assign	vad_gru_input_weights_array[ 1145] = 32'b11000010000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1146] = 32'b01000010111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1147] = 32'b11000010101100100000000000000000;
	assign	vad_gru_input_weights_array[ 1148] = 32'b01000010000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1149] = 32'b11000010110101100000000000000000;
	assign	vad_gru_input_weights_array[ 1150] = 32'b01000010001011000000000000000000;
	assign	vad_gru_input_weights_array[ 1151] = 32'b11000001100010000000000000000000;
	assign	vad_gru_input_weights_array[ 1152] = 32'b01000001110000000000000000000000;
	assign	vad_gru_input_weights_array[ 1153] = 32'b01000001110000000000000000000000;
	assign	vad_gru_input_weights_array[ 1154] = 32'b01000001100100000000000000000000;
	assign	vad_gru_input_weights_array[ 1155] = 32'b01000001111010000000000000000000;
	assign	vad_gru_input_weights_array[ 1156] = 32'b11000001010100000000000000000000;
	assign	vad_gru_input_weights_array[ 1157] = 32'b11000001011100000000000000000000;
	assign	vad_gru_input_weights_array[ 1158] = 32'b11000010000100000000000000000000;
	assign	vad_gru_input_weights_array[ 1159] = 32'b01000010011110000000000000000000;
	assign	vad_gru_input_weights_array[ 1160] = 32'b11000010101101100000000000000000;
	assign	vad_gru_input_weights_array[ 1161] = 32'b01000000100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1162] = 32'b11000010001001000000000000000000;
	assign	vad_gru_input_weights_array[ 1163] = 32'b01000010101111100000000000000000;
	assign	vad_gru_input_weights_array[ 1164] = 32'b01000001111000000000000000000000;
	assign	vad_gru_input_weights_array[ 1165] = 32'b11000001101110000000000000000000;
	assign	vad_gru_input_weights_array[ 1166] = 32'b01000000110000000000000000000000;
	assign	vad_gru_input_weights_array[ 1167] = 32'b01000010001110000000000000000000;
	assign	vad_gru_input_weights_array[ 1168] = 32'b01000010101010000000000000000000;
	assign	vad_gru_input_weights_array[ 1169] = 32'b01000010100001000000000000000000;
	assign	vad_gru_input_weights_array[ 1170] = 32'b01000010100110100000000000000000;
	assign	vad_gru_input_weights_array[ 1171] = 32'b01000010100010000000000000000000;
	assign	vad_gru_input_weights_array[ 1172] = 32'b11000010100011000000000000000000;
	assign	vad_gru_input_weights_array[ 1173] = 32'b10111111100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1174] = 32'b11000001101110000000000000000000;
	assign	vad_gru_input_weights_array[ 1175] = 32'b11000000110000000000000000000000;
	assign	vad_gru_input_weights_array[ 1176] = 32'b01000010100000100000000000000000;
	assign	vad_gru_input_weights_array[ 1177] = 32'b01000010100011000000000000000000;
	assign	vad_gru_input_weights_array[ 1178] = 32'b11000001101010000000000000000000;
	assign	vad_gru_input_weights_array[ 1179] = 32'b01000001000100000000000000000000;
	assign	vad_gru_input_weights_array[ 1180] = 32'b01000010100110100000000000000000;
	assign	vad_gru_input_weights_array[ 1181] = 32'b11000001010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1182] = 32'b01000000000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1183] = 32'b11000010111011000000000000000000;
	assign	vad_gru_input_weights_array[ 1184] = 32'b01000000100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1185] = 32'b01000001000100000000000000000000;
	assign	vad_gru_input_weights_array[ 1186] = 32'b11000010110110000000000000000000;
	assign	vad_gru_input_weights_array[ 1187] = 32'b01000010101010000000000000000000;
	assign	vad_gru_input_weights_array[ 1188] = 32'b01000010010100000000000000000000;
	assign	vad_gru_input_weights_array[ 1189] = 32'b01000000000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1190] = 32'b01000010010100000000000000000000;
	assign	vad_gru_input_weights_array[ 1191] = 32'b01000001010100000000000000000000;
	assign	vad_gru_input_weights_array[ 1192] = 32'b11000001001000000000000000000000;
	assign	vad_gru_input_weights_array[ 1193] = 32'b01000010011010000000000000000000;
	assign	vad_gru_input_weights_array[ 1194] = 32'b11000010110111000000000000000000;
	assign	vad_gru_input_weights_array[ 1195] = 32'b01000001100100000000000000000000;
	assign	vad_gru_input_weights_array[ 1196] = 32'b01000010100001000000000000000000;
	assign	vad_gru_input_weights_array[ 1197] = 32'b11000010101111100000000000000000;
	assign	vad_gru_input_weights_array[ 1198] = 32'b11000001101110000000000000000000;
	assign	vad_gru_input_weights_array[ 1199] = 32'b01000010100011000000000000000000;
	assign	vad_gru_input_weights_array[ 1200] = 32'b01000001111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1201] = 32'b11000000010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1202] = 32'b01000010011000000000000000000000;
	assign	vad_gru_input_weights_array[ 1203] = 32'b01000010011000000000000000000000;
	assign	vad_gru_input_weights_array[ 1204] = 32'b11000000010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1205] = 32'b11000000111000000000000000000000;
	assign	vad_gru_input_weights_array[ 1206] = 32'b00111111100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1207] = 32'b11000001110110000000000000000000;
	assign	vad_gru_input_weights_array[ 1208] = 32'b11000010010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1209] = 32'b11000010011101000000000000000000;
	assign	vad_gru_input_weights_array[ 1210] = 32'b01000010001001000000000000000000;
	assign	vad_gru_input_weights_array[ 1211] = 32'b11000000100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1212] = 32'b01000001001000000000000000000000;
	assign	vad_gru_input_weights_array[ 1213] = 32'b11000010011110000000000000000000;
	assign	vad_gru_input_weights_array[ 1214] = 32'b01000010000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1215] = 32'b11000000111000000000000000000000;
	assign	vad_gru_input_weights_array[ 1216] = 32'b11000001110000000000000000000000;
	assign	vad_gru_input_weights_array[ 1217] = 32'b01000001000100000000000000000000;
	assign	vad_gru_input_weights_array[ 1218] = 32'b11000010010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1219] = 32'b11000010011100000000000000000000;
	assign	vad_gru_input_weights_array[ 1220] = 32'b11000000100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1221] = 32'b01000010100111100000000000000000;
	assign	vad_gru_input_weights_array[ 1222] = 32'b11000001101000000000000000000000;
	assign	vad_gru_input_weights_array[ 1223] = 32'b11000010000110000000000000000000;
	assign	vad_gru_input_weights_array[ 1224] = 32'b11000010100110000000000000000000;
	assign	vad_gru_input_weights_array[ 1225] = 32'b01000010100010000000000000000000;
	assign	vad_gru_input_weights_array[ 1226] = 32'b11000010010001000000000000000000;
	assign	vad_gru_input_weights_array[ 1227] = 32'b11000010110000100000000000000000;
	assign	vad_gru_input_weights_array[ 1228] = 32'b00000000000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1229] = 32'b11000001011100000000000000000000;
	assign	vad_gru_input_weights_array[ 1230] = 32'b01000000101000000000000000000000;
	assign	vad_gru_input_weights_array[ 1231] = 32'b11000010110010000000000000000000;
	assign	vad_gru_input_weights_array[ 1232] = 32'b11000010010001000000000000000000;
	assign	vad_gru_input_weights_array[ 1233] = 32'b11000010101111100000000000000000;
	assign	vad_gru_input_weights_array[ 1234] = 32'b11000010110001100000000000000000;
	assign	vad_gru_input_weights_array[ 1235] = 32'b11000010111001100000000000000000;
	assign	vad_gru_input_weights_array[ 1236] = 32'b11000001000100000000000000000000;
	assign	vad_gru_input_weights_array[ 1237] = 32'b11000010001000000000000000000000;
	assign	vad_gru_input_weights_array[ 1238] = 32'b01000001001000000000000000000000;
	assign	vad_gru_input_weights_array[ 1239] = 32'b01000010110100000000000000000000;
	assign	vad_gru_input_weights_array[ 1240] = 32'b01000001010100000000000000000000;
	assign	vad_gru_input_weights_array[ 1241] = 32'b01000010011000000000000000000000;
	assign	vad_gru_input_weights_array[ 1242] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[ 1243] = 32'b11000001110110000000000000000000;
	assign	vad_gru_input_weights_array[ 1244] = 32'b11000010110110100000000000000000;
	assign	vad_gru_input_weights_array[ 1245] = 32'b11000010101111000000000000000000;
	assign	vad_gru_input_weights_array[ 1246] = 32'b11000010111011000000000000000000;
	assign	vad_gru_input_weights_array[ 1247] = 32'b11000010110011000000000000000000;
	assign	vad_gru_input_weights_array[ 1248] = 32'b11000010001100000000000000000000;
	assign	vad_gru_input_weights_array[ 1249] = 32'b11000010101010100000000000000000;
	assign	vad_gru_input_weights_array[ 1250] = 32'b01000010010100000000000000000000;
	assign	vad_gru_input_weights_array[ 1251] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[ 1252] = 32'b11000000100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1253] = 32'b01000001011000000000000000000000;
	assign	vad_gru_input_weights_array[ 1254] = 32'b01000010011110000000000000000000;
	assign	vad_gru_input_weights_array[ 1255] = 32'b01000010111100100000000000000000;
	assign	vad_gru_input_weights_array[ 1256] = 32'b11000010111101000000000000000000;
	assign	vad_gru_input_weights_array[ 1257] = 32'b11000001110100000000000000000000;
	assign	vad_gru_input_weights_array[ 1258] = 32'b11000010100111100000000000000000;
	assign	vad_gru_input_weights_array[ 1259] = 32'b11000010001010000000000000000000;
	assign	vad_gru_input_weights_array[ 1260] = 32'b11000010000010000000000000000000;
	assign	vad_gru_input_weights_array[ 1261] = 32'b00111111100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1262] = 32'b01000001110010000000000000000000;
	assign	vad_gru_input_weights_array[ 1263] = 32'b11000010000110000000000000000000;
	assign	vad_gru_input_weights_array[ 1264] = 32'b11000010100111100000000000000000;
	assign	vad_gru_input_weights_array[ 1265] = 32'b11000010011010000000000000000000;
	assign	vad_gru_input_weights_array[ 1266] = 32'b11000001111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1267] = 32'b11000001111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1268] = 32'b11000010101101000000000000000000;
	assign	vad_gru_input_weights_array[ 1269] = 32'b11000001111100000000000000000000;
	assign	vad_gru_input_weights_array[ 1270] = 32'b11000010111101100000000000000000;
	assign	vad_gru_input_weights_array[ 1271] = 32'b01000010000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1272] = 32'b11000010011000000000000000000000;
	assign	vad_gru_input_weights_array[ 1273] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1274] = 32'b01000010100001000000000000000000;
	assign	vad_gru_input_weights_array[ 1275] = 32'b01000010111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1276] = 32'b10111111100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1277] = 32'b01000000010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1278] = 32'b01000010101101100000000000000000;
	assign	vad_gru_input_weights_array[ 1279] = 32'b11000010110011100000000000000000;
	assign	vad_gru_input_weights_array[ 1280] = 32'b11000000111000000000000000000000;
	assign	vad_gru_input_weights_array[ 1281] = 32'b01000001101110000000000000000000;
	assign	vad_gru_input_weights_array[ 1282] = 32'b01000010100111000000000000000000;
	assign	vad_gru_input_weights_array[ 1283] = 32'b11000001100100000000000000000000;
	assign	vad_gru_input_weights_array[ 1284] = 32'b01000001000100000000000000000000;
	assign	vad_gru_input_weights_array[ 1285] = 32'b01000010100010100000000000000000;
	assign	vad_gru_input_weights_array[ 1286] = 32'b11000010100010100000000000000000;
	assign	vad_gru_input_weights_array[ 1287] = 32'b01000010100110000000000000000000;
	assign	vad_gru_input_weights_array[ 1288] = 32'b11000010000110000000000000000000;
	assign	vad_gru_input_weights_array[ 1289] = 32'b11000010000001000000000000000000;
	assign	vad_gru_input_weights_array[ 1290] = 32'b11000000000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1291] = 32'b11000010110001000000000000000000;
	assign	vad_gru_input_weights_array[ 1292] = 32'b01000001100100000000000000000000;
	assign	vad_gru_input_weights_array[ 1293] = 32'b01000010110101000000000000000000;
	assign	vad_gru_input_weights_array[ 1294] = 32'b01000010101010000000000000000000;
	assign	vad_gru_input_weights_array[ 1295] = 32'b01000010010111000000000000000000;
	assign	vad_gru_input_weights_array[ 1296] = 32'b01000010101011100000000000000000;
	assign	vad_gru_input_weights_array[ 1297] = 32'b11000010001111000000000000000000;
	assign	vad_gru_input_weights_array[ 1298] = 32'b01000010000011000000000000000000;
	assign	vad_gru_input_weights_array[ 1299] = 32'b11000010111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1300] = 32'b01000010100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1301] = 32'b01000010001001000000000000000000;
	assign	vad_gru_input_weights_array[ 1302] = 32'b11000001011000000000000000000000;
	assign	vad_gru_input_weights_array[ 1303] = 32'b01000010001110000000000000000000;
	assign	vad_gru_input_weights_array[ 1304] = 32'b01000001110010000000000000000000;
	assign	vad_gru_input_weights_array[ 1305] = 32'b11000000000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1306] = 32'b01000010111100000000000000000000;
	assign	vad_gru_input_weights_array[ 1307] = 32'b11000001101010000000000000000000;
	assign	vad_gru_input_weights_array[ 1308] = 32'b01000010101001000000000000000000;
	assign	vad_gru_input_weights_array[ 1309] = 32'b01000001100110000000000000000000;
	assign	vad_gru_input_weights_array[ 1310] = 32'b11000010100111100000000000000000;
	assign	vad_gru_input_weights_array[ 1311] = 32'b11000010000101000000000000000000;
	assign	vad_gru_input_weights_array[ 1312] = 32'b11000000010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1313] = 32'b11000001000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1314] = 32'b11000001100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1315] = 32'b01000001101010000000000000000000;
	assign	vad_gru_input_weights_array[ 1316] = 32'b01000001100110000000000000000000;
	assign	vad_gru_input_weights_array[ 1317] = 32'b11000000101000000000000000000000;
	assign	vad_gru_input_weights_array[ 1318] = 32'b11000001111000000000000000000000;
	assign	vad_gru_input_weights_array[ 1319] = 32'b11000010111000000000000000000000;
	assign	vad_gru_input_weights_array[ 1320] = 32'b01000010000111000000000000000000;
	assign	vad_gru_input_weights_array[ 1321] = 32'b11000000110000000000000000000000;
	assign	vad_gru_input_weights_array[ 1322] = 32'b11000001111100000000000000000000;
	assign	vad_gru_input_weights_array[ 1323] = 32'b01000010010101000000000000000000;
	assign	vad_gru_input_weights_array[ 1324] = 32'b11000010100010100000000000000000;
	assign	vad_gru_input_weights_array[ 1325] = 32'b01000010010101000000000000000000;
	assign	vad_gru_input_weights_array[ 1326] = 32'b01000010001110000000000000000000;
	assign	vad_gru_input_weights_array[ 1327] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[ 1328] = 32'b01000010111101100000000000000000;
	assign	vad_gru_input_weights_array[ 1329] = 32'b01000010100111000000000000000000;
	assign	vad_gru_input_weights_array[ 1330] = 32'b01000001101000000000000000000000;
	assign	vad_gru_input_weights_array[ 1331] = 32'b01000001111000000000000000000000;
	assign	vad_gru_input_weights_array[ 1332] = 32'b11000000111000000000000000000000;
	assign	vad_gru_input_weights_array[ 1333] = 32'b01000010100100100000000000000000;
	assign	vad_gru_input_weights_array[ 1334] = 32'b01000010100100000000000000000000;
	assign	vad_gru_input_weights_array[ 1335] = 32'b01000001100010000000000000000000;
	assign	vad_gru_input_weights_array[ 1336] = 32'b11000010001000000000000000000000;
	assign	vad_gru_input_weights_array[ 1337] = 32'b01000010001001000000000000000000;
	assign	vad_gru_input_weights_array[ 1338] = 32'b01000010110111100000000000000000;
	assign	vad_gru_input_weights_array[ 1339] = 32'b01000010011001000000000000000000;
	assign	vad_gru_input_weights_array[ 1340] = 32'b01000010000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1341] = 32'b11000010101111100000000000000000;
	assign	vad_gru_input_weights_array[ 1342] = 32'b01000001111010000000000000000000;
	assign	vad_gru_input_weights_array[ 1343] = 32'b01000001111000000000000000000000;
	assign	vad_gru_input_weights_array[ 1344] = 32'b11000010000111000000000000000000;
	assign	vad_gru_input_weights_array[ 1345] = 32'b11000010100000100000000000000000;
	assign	vad_gru_input_weights_array[ 1346] = 32'b01000010010110000000000000000000;
	assign	vad_gru_input_weights_array[ 1347] = 32'b11000001101000000000000000000000;
	assign	vad_gru_input_weights_array[ 1348] = 32'b11000010011111000000000000000000;
	assign	vad_gru_input_weights_array[ 1349] = 32'b01000001111010000000000000000000;
	assign	vad_gru_input_weights_array[ 1350] = 32'b11000010100001100000000000000000;
	assign	vad_gru_input_weights_array[ 1351] = 32'b01000000010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1352] = 32'b01000010001100000000000000000000;
	assign	vad_gru_input_weights_array[ 1353] = 32'b11000010011001000000000000000000;
	assign	vad_gru_input_weights_array[ 1354] = 32'b11000010001111000000000000000000;
	assign	vad_gru_input_weights_array[ 1355] = 32'b01000001001100000000000000000000;
	assign	vad_gru_input_weights_array[ 1356] = 32'b01000010011101000000000000000000;
	assign	vad_gru_input_weights_array[ 1357] = 32'b11000001101100000000000000000000;
	assign	vad_gru_input_weights_array[ 1358] = 32'b11000010001100000000000000000000;
	assign	vad_gru_input_weights_array[ 1359] = 32'b01000010011101000000000000000000;
	assign	vad_gru_input_weights_array[ 1360] = 32'b01000010010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1361] = 32'b11000010110010000000000000000000;
	assign	vad_gru_input_weights_array[ 1362] = 32'b01000001101000000000000000000000;
	assign	vad_gru_input_weights_array[ 1363] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1364] = 32'b01000010110000000000000000000000;
	assign	vad_gru_input_weights_array[ 1365] = 32'b11000001110000000000000000000000;
	assign	vad_gru_input_weights_array[ 1366] = 32'b11000001100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1367] = 32'b01000000010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1368] = 32'b11000010100010100000000000000000;
	assign	vad_gru_input_weights_array[ 1369] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[ 1370] = 32'b01000010100101000000000000000000;
	assign	vad_gru_input_weights_array[ 1371] = 32'b11000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1372] = 32'b01000001000100000000000000000000;
	assign	vad_gru_input_weights_array[ 1373] = 32'b01000010001101000000000000000000;
	assign	vad_gru_input_weights_array[ 1374] = 32'b11000010100001100000000000000000;
	assign	vad_gru_input_weights_array[ 1375] = 32'b11000010111101100000000000000000;
	assign	vad_gru_input_weights_array[ 1376] = 32'b11000010011011000000000000000000;
	assign	vad_gru_input_weights_array[ 1377] = 32'b11000010100100000000000000000000;
	assign	vad_gru_input_weights_array[ 1378] = 32'b01000010111011000000000000000000;
	assign	vad_gru_input_weights_array[ 1379] = 32'b01000010100010100000000000000000;
	assign	vad_gru_input_weights_array[ 1380] = 32'b01000010001101000000000000000000;
	assign	vad_gru_input_weights_array[ 1381] = 32'b01000010010010000000000000000000;
	assign	vad_gru_input_weights_array[ 1382] = 32'b11000010011001000000000000000000;
	assign	vad_gru_input_weights_array[ 1383] = 32'b01000010100001100000000000000000;
	assign	vad_gru_input_weights_array[ 1384] = 32'b01000001010100000000000000000000;
	assign	vad_gru_input_weights_array[ 1385] = 32'b11000010100001000000000000000000;
	assign	vad_gru_input_weights_array[ 1386] = 32'b11000010110101000000000000000000;
	assign	vad_gru_input_weights_array[ 1387] = 32'b01000010001111000000000000000000;
	assign	vad_gru_input_weights_array[ 1388] = 32'b01000010011110000000000000000000;
	assign	vad_gru_input_weights_array[ 1389] = 32'b01000001101100000000000000000000;
	assign	vad_gru_input_weights_array[ 1390] = 32'b10111111100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1391] = 32'b11000001101100000000000000000000;
	assign	vad_gru_input_weights_array[ 1392] = 32'b11000001110010000000000000000000;
	assign	vad_gru_input_weights_array[ 1393] = 32'b11000010001000000000000000000000;
	assign	vad_gru_input_weights_array[ 1394] = 32'b11000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1395] = 32'b01000000010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1396] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1397] = 32'b01000010000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1398] = 32'b01000010110011000000000000000000;
	assign	vad_gru_input_weights_array[ 1399] = 32'b11000010011000000000000000000000;
	assign	vad_gru_input_weights_array[ 1400] = 32'b11000001110010000000000000000000;
	assign	vad_gru_input_weights_array[ 1401] = 32'b11000010100101100000000000000000;
	assign	vad_gru_input_weights_array[ 1402] = 32'b11000001111100000000000000000000;
	assign	vad_gru_input_weights_array[ 1403] = 32'b01000010111101000000000000000000;
	assign	vad_gru_input_weights_array[ 1404] = 32'b01000010011100000000000000000000;
	assign	vad_gru_input_weights_array[ 1405] = 32'b11000001010100000000000000000000;
	assign	vad_gru_input_weights_array[ 1406] = 32'b01000010000100000000000000000000;
	assign	vad_gru_input_weights_array[ 1407] = 32'b11000010100100100000000000000000;
	assign	vad_gru_input_weights_array[ 1408] = 32'b01000000111000000000000000000000;
	assign	vad_gru_input_weights_array[ 1409] = 32'b11000010101010000000000000000000;
	assign	vad_gru_input_weights_array[ 1410] = 32'b01000010111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1411] = 32'b01000010001000000000000000000000;
	assign	vad_gru_input_weights_array[ 1412] = 32'b11000010111011000000000000000000;
	assign	vad_gru_input_weights_array[ 1413] = 32'b01000001100010000000000000000000;
	assign	vad_gru_input_weights_array[ 1414] = 32'b11000010101011100000000000000000;
	assign	vad_gru_input_weights_array[ 1415] = 32'b11000010111011000000000000000000;
	assign	vad_gru_input_weights_array[ 1416] = 32'b11000001000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1417] = 32'b01000000010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1418] = 32'b11000001110110000000000000000000;
	assign	vad_gru_input_weights_array[ 1419] = 32'b01000010110111100000000000000000;
	assign	vad_gru_input_weights_array[ 1420] = 32'b11000010001000000000000000000000;
	assign	vad_gru_input_weights_array[ 1421] = 32'b01000010001000000000000000000000;
	assign	vad_gru_input_weights_array[ 1422] = 32'b11000010010011000000000000000000;
	assign	vad_gru_input_weights_array[ 1423] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[ 1424] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1425] = 32'b11000010001101000000000000000000;
	assign	vad_gru_input_weights_array[ 1426] = 32'b11000001111100000000000000000000;
	assign	vad_gru_input_weights_array[ 1427] = 32'b11000010010110000000000000000000;
	assign	vad_gru_input_weights_array[ 1428] = 32'b01000010001110000000000000000000;
	assign	vad_gru_input_weights_array[ 1429] = 32'b01000010101000000000000000000000;
	assign	vad_gru_input_weights_array[ 1430] = 32'b10111111100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1431] = 32'b11000001111100000000000000000000;
	assign	vad_gru_input_weights_array[ 1432] = 32'b01000010110010100000000000000000;
	assign	vad_gru_input_weights_array[ 1433] = 32'b11000001100010000000000000000000;
	assign	vad_gru_input_weights_array[ 1434] = 32'b01000001100100000000000000000000;
	assign	vad_gru_input_weights_array[ 1435] = 32'b01000001110100000000000000000000;
	assign	vad_gru_input_weights_array[ 1436] = 32'b01000010010110000000000000000000;
	assign	vad_gru_input_weights_array[ 1437] = 32'b01000000111000000000000000000000;
	assign	vad_gru_input_weights_array[ 1438] = 32'b11000001010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1439] = 32'b00111111100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1440] = 32'b11000010111111100000000000000000;
	assign	vad_gru_input_weights_array[ 1441] = 32'b01000010111101100000000000000000;
	assign	vad_gru_input_weights_array[ 1442] = 32'b11000010111101000000000000000000;
	assign	vad_gru_input_weights_array[ 1443] = 32'b11000001110110000000000000000000;
	assign	vad_gru_input_weights_array[ 1444] = 32'b11000010100101100000000000000000;
	assign	vad_gru_input_weights_array[ 1445] = 32'b01000010100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1446] = 32'b01000001001000000000000000000000;
	assign	vad_gru_input_weights_array[ 1447] = 32'b01000001110010000000000000000000;
	assign	vad_gru_input_weights_array[ 1448] = 32'b11000001011100000000000000000000;
	assign	vad_gru_input_weights_array[ 1449] = 32'b11000010001100000000000000000000;
	assign	vad_gru_input_weights_array[ 1450] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[ 1451] = 32'b11000010111111100000000000000000;
	assign	vad_gru_input_weights_array[ 1452] = 32'b01000000101000000000000000000000;
	assign	vad_gru_input_weights_array[ 1453] = 32'b11000010101010000000000000000000;
	assign	vad_gru_input_weights_array[ 1454] = 32'b11000010101000100000000000000000;
	assign	vad_gru_input_weights_array[ 1455] = 32'b11000000111000000000000000000000;
	assign	vad_gru_input_weights_array[ 1456] = 32'b01000001100110000000000000000000;
	assign	vad_gru_input_weights_array[ 1457] = 32'b11000001110100000000000000000000;
	assign	vad_gru_input_weights_array[ 1458] = 32'b01000010111111000000000000000000;
	assign	vad_gru_input_weights_array[ 1459] = 32'b01000001011100000000000000000000;
	assign	vad_gru_input_weights_array[ 1460] = 32'b01000010111010000000000000000000;
	assign	vad_gru_input_weights_array[ 1461] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[ 1462] = 32'b01000001011000000000000000000000;
	assign	vad_gru_input_weights_array[ 1463] = 32'b11000010100110000000000000000000;
	assign	vad_gru_input_weights_array[ 1464] = 32'b01000010001100000000000000000000;
	assign	vad_gru_input_weights_array[ 1465] = 32'b01000010011110000000000000000000;
	assign	vad_gru_input_weights_array[ 1466] = 32'b11000010110111000000000000000000;
	assign	vad_gru_input_weights_array[ 1467] = 32'b11000010111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1468] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1469] = 32'b11000001111010000000000000000000;
	assign	vad_gru_input_weights_array[ 1470] = 32'b11000010101011100000000000000000;
	assign	vad_gru_input_weights_array[ 1471] = 32'b11000000010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1472] = 32'b11000010100010100000000000000000;
	assign	vad_gru_input_weights_array[ 1473] = 32'b01000010101001000000000000000000;
	assign	vad_gru_input_weights_array[ 1474] = 32'b01000010101101000000000000000000;
	assign	vad_gru_input_weights_array[ 1475] = 32'b01000010011001000000000000000000;
	assign	vad_gru_input_weights_array[ 1476] = 32'b11000010111101100000000000000000;
	assign	vad_gru_input_weights_array[ 1477] = 32'b01000010111101100000000000000000;
	assign	vad_gru_input_weights_array[ 1478] = 32'b01000010110010000000000000000000;
	assign	vad_gru_input_weights_array[ 1479] = 32'b11000001100110000000000000000000;
	assign	vad_gru_input_weights_array[ 1480] = 32'b11000010010011000000000000000000;
	assign	vad_gru_input_weights_array[ 1481] = 32'b11000010000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1482] = 32'b01000010100010100000000000000000;
	assign	vad_gru_input_weights_array[ 1483] = 32'b01000010000101000000000000000000;
	assign	vad_gru_input_weights_array[ 1484] = 32'b11000010011001000000000000000000;
	assign	vad_gru_input_weights_array[ 1485] = 32'b11000011000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1486] = 32'b11000010111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1487] = 32'b11000010100100000000000000000000;
	assign	vad_gru_input_weights_array[ 1488] = 32'b11000001010100000000000000000000;
	assign	vad_gru_input_weights_array[ 1489] = 32'b01000010010011000000000000000000;
	assign	vad_gru_input_weights_array[ 1490] = 32'b11000000111000000000000000000000;
	assign	vad_gru_input_weights_array[ 1491] = 32'b11000010001101000000000000000000;
	assign	vad_gru_input_weights_array[ 1492] = 32'b11000010100100100000000000000000;
	assign	vad_gru_input_weights_array[ 1493] = 32'b01000000101000000000000000000000;
	assign	vad_gru_input_weights_array[ 1494] = 32'b01000010110001100000000000000000;
	assign	vad_gru_input_weights_array[ 1495] = 32'b11000001110100000000000000000000;
	assign	vad_gru_input_weights_array[ 1496] = 32'b11000010111010100000000000000000;
	assign	vad_gru_input_weights_array[ 1497] = 32'b11000010110000000000000000000000;
	assign	vad_gru_input_weights_array[ 1498] = 32'b11000010110110100000000000000000;
	assign	vad_gru_input_weights_array[ 1499] = 32'b01000000100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1500] = 32'b11000001111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1501] = 32'b11000001010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1502] = 32'b00000000000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1503] = 32'b01000001111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1504] = 32'b11000010001010000000000000000000;
	assign	vad_gru_input_weights_array[ 1505] = 32'b11000001110110000000000000000000;
	assign	vad_gru_input_weights_array[ 1506] = 32'b01000001010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1507] = 32'b11000010101000100000000000000000;
	assign	vad_gru_input_weights_array[ 1508] = 32'b01000010111011000000000000000000;
	assign	vad_gru_input_weights_array[ 1509] = 32'b01000010000111000000000000000000;
	assign	vad_gru_input_weights_array[ 1510] = 32'b01000010101001100000000000000000;
	assign	vad_gru_input_weights_array[ 1511] = 32'b01000001011000000000000000000000;
	assign	vad_gru_input_weights_array[ 1512] = 32'b01000010001001000000000000000000;
	assign	vad_gru_input_weights_array[ 1513] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[ 1514] = 32'b01000010110101100000000000000000;
	assign	vad_gru_input_weights_array[ 1515] = 32'b11000010101001000000000000000000;
	assign	vad_gru_input_weights_array[ 1516] = 32'b01000010101111000000000000000000;
	assign	vad_gru_input_weights_array[ 1517] = 32'b11000010111010000000000000000000;
	assign	vad_gru_input_weights_array[ 1518] = 32'b11000010111101000000000000000000;
	assign	vad_gru_input_weights_array[ 1519] = 32'b11000010001111000000000000000000;
	assign	vad_gru_input_weights_array[ 1520] = 32'b11000010110110100000000000000000;
	assign	vad_gru_input_weights_array[ 1521] = 32'b11000010101010000000000000000000;
	assign	vad_gru_input_weights_array[ 1522] = 32'b11000011000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1523] = 32'b11000010000011000000000000000000;
	assign	vad_gru_input_weights_array[ 1524] = 32'b11000010011000000000000000000000;
	assign	vad_gru_input_weights_array[ 1525] = 32'b01000010100001000000000000000000;
	assign	vad_gru_input_weights_array[ 1526] = 32'b01000001000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1527] = 32'b11000010100000100000000000000000;
	assign	vad_gru_input_weights_array[ 1528] = 32'b01000001100110000000000000000000;
	assign	vad_gru_input_weights_array[ 1529] = 32'b01000010001010000000000000000000;
	assign	vad_gru_input_weights_array[ 1530] = 32'b11000010001110000000000000000000;
	assign	vad_gru_input_weights_array[ 1531] = 32'b11000010100100000000000000000000;
	assign	vad_gru_input_weights_array[ 1532] = 32'b11000010110110100000000000000000;
	assign	vad_gru_input_weights_array[ 1533] = 32'b01000010001001000000000000000000;
	assign	vad_gru_input_weights_array[ 1534] = 32'b01000010001011000000000000000000;
	assign	vad_gru_input_weights_array[ 1535] = 32'b11000010111111100000000000000000;
	assign	vad_gru_input_weights_array[ 1536] = 32'b11000010111000100000000000000000;
	assign	vad_gru_input_weights_array[ 1537] = 32'b01000010011010000000000000000000;
	assign	vad_gru_input_weights_array[ 1538] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[ 1539] = 32'b01000010001010000000000000000000;
	assign	vad_gru_input_weights_array[ 1540] = 32'b11000010100101100000000000000000;
	assign	vad_gru_input_weights_array[ 1541] = 32'b10111111100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1542] = 32'b01000010100000100000000000000000;
	assign	vad_gru_input_weights_array[ 1543] = 32'b01000010111010100000000000000000;
	assign	vad_gru_input_weights_array[ 1544] = 32'b11000010010111000000000000000000;
	assign	vad_gru_input_weights_array[ 1545] = 32'b11000010111000100000000000000000;
	assign	vad_gru_input_weights_array[ 1546] = 32'b11000010111101100000000000000000;
	assign	vad_gru_input_weights_array[ 1547] = 32'b01000010111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1548] = 32'b01000010001011000000000000000000;
	assign	vad_gru_input_weights_array[ 1549] = 32'b11000010110000000000000000000000;
	assign	vad_gru_input_weights_array[ 1550] = 32'b11000010111001100000000000000000;
	assign	vad_gru_input_weights_array[ 1551] = 32'b11000001100110000000000000000000;
	assign	vad_gru_input_weights_array[ 1552] = 32'b01000010100010000000000000000000;
	assign	vad_gru_input_weights_array[ 1553] = 32'b01000001011100000000000000000000;
	assign	vad_gru_input_weights_array[ 1554] = 32'b01000010101111000000000000000000;
	assign	vad_gru_input_weights_array[ 1555] = 32'b01000000010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1556] = 32'b01000010100101100000000000000000;
	assign	vad_gru_input_weights_array[ 1557] = 32'b00000000000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1558] = 32'b01000010000010000000000000000000;
	assign	vad_gru_input_weights_array[ 1559] = 32'b01000001000100000000000000000000;
	assign	vad_gru_input_weights_array[ 1560] = 32'b01000010001010000000000000000000;
	assign	vad_gru_input_weights_array[ 1561] = 32'b01000010110111000000000000000000;
	assign	vad_gru_input_weights_array[ 1562] = 32'b11000010010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1563] = 32'b01000010101110000000000000000000;
	assign	vad_gru_input_weights_array[ 1564] = 32'b11000010100110000000000000000000;
	assign	vad_gru_input_weights_array[ 1565] = 32'b01000010110001100000000000000000;
	assign	vad_gru_input_weights_array[ 1566] = 32'b11000001100010000000000000000000;
	assign	vad_gru_input_weights_array[ 1567] = 32'b01000001110110000000000000000000;
	assign	vad_gru_input_weights_array[ 1568] = 32'b01000010000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1569] = 32'b01000001010100000000000000000000;
	assign	vad_gru_input_weights_array[ 1570] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1571] = 32'b01000010010010000000000000000000;
	assign	vad_gru_input_weights_array[ 1572] = 32'b11000001100010000000000000000000;
	assign	vad_gru_input_weights_array[ 1573] = 32'b01000010011000000000000000000000;
	assign	vad_gru_input_weights_array[ 1574] = 32'b01000000100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1575] = 32'b01000010010101000000000000000000;
	assign	vad_gru_input_weights_array[ 1576] = 32'b01000010000010000000000000000000;
	assign	vad_gru_input_weights_array[ 1577] = 32'b11000001000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1578] = 32'b01000010110001100000000000000000;
	assign	vad_gru_input_weights_array[ 1579] = 32'b01000010101000000000000000000000;
	assign	vad_gru_input_weights_array[ 1580] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[ 1581] = 32'b11000001101010000000000000000000;
	assign	vad_gru_input_weights_array[ 1582] = 32'b11000010100000100000000000000000;
	assign	vad_gru_input_weights_array[ 1583] = 32'b11000001001100000000000000000000;
	assign	vad_gru_input_weights_array[ 1584] = 32'b11000010001110000000000000000000;
	assign	vad_gru_input_weights_array[ 1585] = 32'b01000010001100000000000000000000;
	assign	vad_gru_input_weights_array[ 1586] = 32'b11000010101000100000000000000000;
	assign	vad_gru_input_weights_array[ 1587] = 32'b11000000010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1588] = 32'b11000010111100100000000000000000;
	assign	vad_gru_input_weights_array[ 1589] = 32'b01000010111101100000000000000000;
	assign	vad_gru_input_weights_array[ 1590] = 32'b01000010100001000000000000000000;
	assign	vad_gru_input_weights_array[ 1591] = 32'b11000010101000100000000000000000;
	assign	vad_gru_input_weights_array[ 1592] = 32'b11000010101010000000000000000000;
	assign	vad_gru_input_weights_array[ 1593] = 32'b01000010111011100000000000000000;
	assign	vad_gru_input_weights_array[ 1594] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[ 1595] = 32'b01000010101010000000000000000000;
	assign	vad_gru_input_weights_array[ 1596] = 32'b01000010110100100000000000000000;
	assign	vad_gru_input_weights_array[ 1597] = 32'b01000010001101000000000000000000;
	assign	vad_gru_input_weights_array[ 1598] = 32'b11000010100001000000000000000000;
	assign	vad_gru_input_weights_array[ 1599] = 32'b11000010001010000000000000000000;
	assign	vad_gru_input_weights_array[ 1600] = 32'b11000001101110000000000000000000;
	assign	vad_gru_input_weights_array[ 1601] = 32'b01000010000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1602] = 32'b11000001110010000000000000000000;
	assign	vad_gru_input_weights_array[ 1603] = 32'b01000001010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1604] = 32'b01000010110111100000000000000000;
	assign	vad_gru_input_weights_array[ 1605] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[ 1606] = 32'b01000010101100000000000000000000;
	assign	vad_gru_input_weights_array[ 1607] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1608] = 32'b01000001111100000000000000000000;
	assign	vad_gru_input_weights_array[ 1609] = 32'b01000001110000000000000000000000;
	assign	vad_gru_input_weights_array[ 1610] = 32'b11000010111111100000000000000000;
	assign	vad_gru_input_weights_array[ 1611] = 32'b11000001000100000000000000000000;
	assign	vad_gru_input_weights_array[ 1612] = 32'b11000010010110000000000000000000;
	assign	vad_gru_input_weights_array[ 1613] = 32'b01000010111111100000000000000000;
	assign	vad_gru_input_weights_array[ 1614] = 32'b11000010111010000000000000000000;
	assign	vad_gru_input_weights_array[ 1615] = 32'b11000010111011100000000000000000;
	assign	vad_gru_input_weights_array[ 1616] = 32'b01000010101100000000000000000000;
	assign	vad_gru_input_weights_array[ 1617] = 32'b01000010100011000000000000000000;
	assign	vad_gru_input_weights_array[ 1618] = 32'b01000010101111000000000000000000;
	assign	vad_gru_input_weights_array[ 1619] = 32'b11000010111100000000000000000000;
	assign	vad_gru_input_weights_array[ 1620] = 32'b01000010000011000000000000000000;
	assign	vad_gru_input_weights_array[ 1621] = 32'b11000010101110100000000000000000;
	assign	vad_gru_input_weights_array[ 1622] = 32'b01000001011100000000000000000000;
	assign	vad_gru_input_weights_array[ 1623] = 32'b01000001101100000000000000000000;
	assign	vad_gru_input_weights_array[ 1624] = 32'b11000001101010000000000000000000;
	assign	vad_gru_input_weights_array[ 1625] = 32'b01000001110010000000000000000000;
	assign	vad_gru_input_weights_array[ 1626] = 32'b11000010110111000000000000000000;
	assign	vad_gru_input_weights_array[ 1627] = 32'b11000010111101100000000000000000;
	assign	vad_gru_input_weights_array[ 1628] = 32'b11000010001101000000000000000000;
	assign	vad_gru_input_weights_array[ 1629] = 32'b01000001000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1630] = 32'b11000010110110100000000000000000;
	assign	vad_gru_input_weights_array[ 1631] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1632] = 32'b11000010111101000000000000000000;
	assign	vad_gru_input_weights_array[ 1633] = 32'b11000010101011000000000000000000;
	assign	vad_gru_input_weights_array[ 1634] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[ 1635] = 32'b01000001000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1636] = 32'b11000001011000000000000000000000;
	assign	vad_gru_input_weights_array[ 1637] = 32'b11000010111100000000000000000000;
	assign	vad_gru_input_weights_array[ 1638] = 32'b11000010001101000000000000000000;
	assign	vad_gru_input_weights_array[ 1639] = 32'b11000010001101000000000000000000;
	assign	vad_gru_input_weights_array[ 1640] = 32'b01000010100010100000000000000000;
	assign	vad_gru_input_weights_array[ 1641] = 32'b11000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1642] = 32'b11000010111101000000000000000000;
	assign	vad_gru_input_weights_array[ 1643] = 32'b01000000110000000000000000000000;
	assign	vad_gru_input_weights_array[ 1644] = 32'b01000010101000100000000000000000;
	assign	vad_gru_input_weights_array[ 1645] = 32'b01000010101011000000000000000000;
	assign	vad_gru_input_weights_array[ 1646] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1647] = 32'b01000010101111100000000000000000;
	assign	vad_gru_input_weights_array[ 1648] = 32'b01000010010110000000000000000000;
	assign	vad_gru_input_weights_array[ 1649] = 32'b01000010100110100000000000000000;
	assign	vad_gru_input_weights_array[ 1650] = 32'b01000010010110000000000000000000;
	assign	vad_gru_input_weights_array[ 1651] = 32'b11000010111101100000000000000000;
	assign	vad_gru_input_weights_array[ 1652] = 32'b01000010111111000000000000000000;
	assign	vad_gru_input_weights_array[ 1653] = 32'b11000010101010100000000000000000;
	assign	vad_gru_input_weights_array[ 1654] = 32'b11000010111010100000000000000000;
	assign	vad_gru_input_weights_array[ 1655] = 32'b01000010011000000000000000000000;
	assign	vad_gru_input_weights_array[ 1656] = 32'b01000001001100000000000000000000;
	assign	vad_gru_input_weights_array[ 1657] = 32'b00000000000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1658] = 32'b11000010011101000000000000000000;
	assign	vad_gru_input_weights_array[ 1659] = 32'b11000010101101100000000000000000;
	assign	vad_gru_input_weights_array[ 1660] = 32'b11000001010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1661] = 32'b11000000000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1662] = 32'b11000010111000100000000000000000;
	assign	vad_gru_input_weights_array[ 1663] = 32'b11000000010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1664] = 32'b11000001011100000000000000000000;
	assign	vad_gru_input_weights_array[ 1665] = 32'b11000010111101000000000000000000;
	assign	vad_gru_input_weights_array[ 1666] = 32'b11000010011111000000000000000000;
	assign	vad_gru_input_weights_array[ 1667] = 32'b11000010101101100000000000000000;
	assign	vad_gru_input_weights_array[ 1668] = 32'b01000001001000000000000000000000;
	assign	vad_gru_input_weights_array[ 1669] = 32'b01000010101010000000000000000000;
	assign	vad_gru_input_weights_array[ 1670] = 32'b11000010110111100000000000000000;
	assign	vad_gru_input_weights_array[ 1671] = 32'b01000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1672] = 32'b01000010101110100000000000000000;
	assign	vad_gru_input_weights_array[ 1673] = 32'b01000001101010000000000000000000;
	assign	vad_gru_input_weights_array[ 1674] = 32'b01000010011110000000000000000000;
	assign	vad_gru_input_weights_array[ 1675] = 32'b11000010100111000000000000000000;
	assign	vad_gru_input_weights_array[ 1676] = 32'b11000010111010000000000000000000;
	assign	vad_gru_input_weights_array[ 1677] = 32'b01000001010100000000000000000000;
	assign	vad_gru_input_weights_array[ 1678] = 32'b11000010011001000000000000000000;
	assign	vad_gru_input_weights_array[ 1679] = 32'b01000001111000000000000000000000;
	assign	vad_gru_input_weights_array[ 1680] = 32'b11000010111110000000000000000000;
	assign	vad_gru_input_weights_array[ 1681] = 32'b01000010111111000000000000000000;
	assign	vad_gru_input_weights_array[ 1682] = 32'b01000010110111000000000000000000;
	assign	vad_gru_input_weights_array[ 1683] = 32'b01000001010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1684] = 32'b01000001011100000000000000000000;
	assign	vad_gru_input_weights_array[ 1685] = 32'b01000010101111100000000000000000;
	assign	vad_gru_input_weights_array[ 1686] = 32'b01000001011100000000000000000000;
	assign	vad_gru_input_weights_array[ 1687] = 32'b11000001100110000000000000000000;
	assign	vad_gru_input_weights_array[ 1688] = 32'b11000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1689] = 32'b11000010110000100000000000000000;
	assign	vad_gru_input_weights_array[ 1690] = 32'b01000010010100000000000000000000;
	assign	vad_gru_input_weights_array[ 1691] = 32'b11000000111000000000000000000000;
	assign	vad_gru_input_weights_array[ 1692] = 32'b01000010110010100000000000000000;
	assign	vad_gru_input_weights_array[ 1693] = 32'b01000001000100000000000000000000;
	assign	vad_gru_input_weights_array[ 1694] = 32'b01000001101000000000000000000000;
	assign	vad_gru_input_weights_array[ 1695] = 32'b11000010111110100000000000000000;
	assign	vad_gru_input_weights_array[ 1696] = 32'b11000001110100000000000000000000;
	assign	vad_gru_input_weights_array[ 1697] = 32'b11000010011000000000000000000000;
	assign	vad_gru_input_weights_array[ 1698] = 32'b01000010100100000000000000000000;
	assign	vad_gru_input_weights_array[ 1699] = 32'b01000010100110100000000000000000;
	assign	vad_gru_input_weights_array[ 1700] = 32'b01000001010000000000000000000000;
	assign	vad_gru_input_weights_array[ 1701] = 32'b11000010111111000000000000000000;
	assign	vad_gru_input_weights_array[ 1702] = 32'b01000001101100000000000000000000;
	assign	vad_gru_input_weights_array[ 1703] = 32'b11000001111010000000000000000000;
	assign	vad_gru_input_weights_array[ 1704] = 32'b01000010001111000000000000000000;
	assign	vad_gru_input_weights_array[ 1705] = 32'b01000010011110000000000000000000;
	assign	vad_gru_input_weights_array[ 1706] = 32'b01000010101111100000000000000000;
	assign	vad_gru_input_weights_array[ 1707] = 32'b01000010111000000000000000000000;
	assign	vad_gru_input_weights_array[ 1708] = 32'b01000010100010100000000000000000;
	assign	vad_gru_input_weights_array[ 1709] = 32'b01000010000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1710] = 32'b01000010110000100000000000000000;
	assign	vad_gru_input_weights_array[ 1711] = 32'b11000010101001100000000000000000;
	assign	vad_gru_input_weights_array[ 1712] = 32'b11000001000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1713] = 32'b11000000101000000000000000000000;
	assign	vad_gru_input_weights_array[ 1714] = 32'b01000010100001100000000000000000;
	assign	vad_gru_input_weights_array[ 1715] = 32'b11000010011111000000000000000000;
	assign	vad_gru_input_weights_array[ 1716] = 32'b11000010111101100000000000000000;
	assign	vad_gru_input_weights_array[ 1717] = 32'b01000010100111100000000000000000;
	assign	vad_gru_input_weights_array[ 1718] = 32'b01000010011011000000000000000000;
	assign	vad_gru_input_weights_array[ 1719] = 32'b00000000000000000000000000000000;
	assign	vad_gru_input_weights_array[ 1720] = 32'b11000000110000000000000000000000;
	assign	vad_gru_input_weights_array[ 1721] = 32'b11000001100010000000000000000000;
	assign	vad_gru_input_weights_array[ 1722] = 32'b01000000100000000000000000000000;
	assign	vad_gru_input_weights_array[ 1723] = 32'b11000010110111100000000000000000;
	assign	vad_gru_input_weights_array[ 1724] = 32'b11000010010100000000000000000000;
	assign	vad_gru_input_weights_array[ 1725] = 32'b01000001110110000000000000000000;
	assign	vad_gru_input_weights_array[ 1726] = 32'b01000010100000100000000000000000;
	assign	vad_gru_input_weights_array[ 1727] = 32'b00000000000000000000000000000000;

	assign	vad_gru_recurrent_weights_array[    0] = 32'b01000010100000100000000000000000;
	assign	vad_gru_recurrent_weights_array[    1] = 32'b01000010101001100000000000000000;
	assign	vad_gru_recurrent_weights_array[    2] = 32'b01000010000011000000000000000000;
	assign	vad_gru_recurrent_weights_array[    3] = 32'b01000010011000000000000000000000;
	assign	vad_gru_recurrent_weights_array[    4] = 32'b01000001110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[    5] = 32'b11000010000010000000000000000000;
	assign	vad_gru_recurrent_weights_array[    6] = 32'b11000001111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[    7] = 32'b11000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[    8] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[    9] = 32'b01000001100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[   10] = 32'b01000010001010000000000000000000;
	assign	vad_gru_recurrent_weights_array[   11] = 32'b11000001000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[   12] = 32'b01000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[   13] = 32'b11000010010101000000000000000000;
	assign	vad_gru_recurrent_weights_array[   14] = 32'b01000001110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[   15] = 32'b11000010101011100000000000000000;
	assign	vad_gru_recurrent_weights_array[   16] = 32'b01000001001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[   17] = 32'b01000010000011000000000000000000;
	assign	vad_gru_recurrent_weights_array[   18] = 32'b11000010101000100000000000000000;
	assign	vad_gru_recurrent_weights_array[   19] = 32'b11000010000011000000000000000000;
	assign	vad_gru_recurrent_weights_array[   20] = 32'b11000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[   21] = 32'b11000001111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[   22] = 32'b01000010111101100000000000000000;
	assign	vad_gru_recurrent_weights_array[   23] = 32'b11000001101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[   24] = 32'b01000010000001000000000000000000;
	assign	vad_gru_recurrent_weights_array[   25] = 32'b11000010101101100000000000000000;
	assign	vad_gru_recurrent_weights_array[   26] = 32'b01000010111000100000000000000000;
	assign	vad_gru_recurrent_weights_array[   27] = 32'b11000010101110100000000000000000;
	assign	vad_gru_recurrent_weights_array[   28] = 32'b01000010001101000000000000000000;
	assign	vad_gru_recurrent_weights_array[   29] = 32'b11000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[   30] = 32'b01000010010101000000000000000000;
	assign	vad_gru_recurrent_weights_array[   31] = 32'b01000010000110000000000000000000;
	assign	vad_gru_recurrent_weights_array[   32] = 32'b11000010101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[   33] = 32'b01000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[   34] = 32'b11000001110110000000000000000000;
	assign	vad_gru_recurrent_weights_array[   35] = 32'b01000010101011100000000000000000;
	assign	vad_gru_recurrent_weights_array[   36] = 32'b01000000100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[   37] = 32'b01000010001011000000000000000000;
	assign	vad_gru_recurrent_weights_array[   38] = 32'b01000010001011000000000000000000;
	assign	vad_gru_recurrent_weights_array[   39] = 32'b01000001001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[   40] = 32'b11000011000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[   41] = 32'b11000011000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[   42] = 32'b11000010001110000000000000000000;
	assign	vad_gru_recurrent_weights_array[   43] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[   44] = 32'b11000010000110000000000000000000;
	assign	vad_gru_recurrent_weights_array[   45] = 32'b11000010001101000000000000000000;
	assign	vad_gru_recurrent_weights_array[   46] = 32'b01000001110010000000000000000000;
	assign	vad_gru_recurrent_weights_array[   47] = 32'b11000010101011100000000000000000;
	assign	vad_gru_recurrent_weights_array[   48] = 32'b01000001100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[   49] = 32'b01000000101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[   50] = 32'b01000010010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[   51] = 32'b11000010110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[   52] = 32'b11000001101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[   53] = 32'b11000001111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[   54] = 32'b01000010111100100000000000000000;
	assign	vad_gru_recurrent_weights_array[   55] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[   56] = 32'b11000001110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[   57] = 32'b11000001101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[   58] = 32'b11000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[   59] = 32'b01000010100010100000000000000000;
	assign	vad_gru_recurrent_weights_array[   60] = 32'b11000010010010000000000000000000;
	assign	vad_gru_recurrent_weights_array[   61] = 32'b01000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[   62] = 32'b01000010100011100000000000000000;
	assign	vad_gru_recurrent_weights_array[   63] = 32'b11000010101000100000000000000000;
	assign	vad_gru_recurrent_weights_array[   64] = 32'b11000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[   65] = 32'b01000010101101000000000000000000;
	assign	vad_gru_recurrent_weights_array[   66] = 32'b11000010101111000000000000000000;
	assign	vad_gru_recurrent_weights_array[   67] = 32'b00111111100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[   68] = 32'b11000010000110000000000000000000;
	assign	vad_gru_recurrent_weights_array[   69] = 32'b01000010000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[   70] = 32'b01000010101100100000000000000000;
	assign	vad_gru_recurrent_weights_array[   71] = 32'b01000001100010000000000000000000;
	assign	vad_gru_recurrent_weights_array[   72] = 32'b11000010011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[   73] = 32'b01000010100011100000000000000000;
	assign	vad_gru_recurrent_weights_array[   74] = 32'b11000010010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[   75] = 32'b01000001100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[   76] = 32'b11000001011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[   77] = 32'b01000010001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[   78] = 32'b11000001100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[   79] = 32'b01000010011011000000000000000000;
	assign	vad_gru_recurrent_weights_array[   80] = 32'b01000001001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[   81] = 32'b01000010111001000000000000000000;
	assign	vad_gru_recurrent_weights_array[   82] = 32'b11000010010011000000000000000000;
	assign	vad_gru_recurrent_weights_array[   83] = 32'b01000010000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[   84] = 32'b01000010110111000000000000000000;
	assign	vad_gru_recurrent_weights_array[   85] = 32'b00111111100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[   86] = 32'b01000000100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[   87] = 32'b01000010110110100000000000000000;
	assign	vad_gru_recurrent_weights_array[   88] = 32'b11000001110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[   89] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[   90] = 32'b01000001110110000000000000000000;
	assign	vad_gru_recurrent_weights_array[   91] = 32'b01000010011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[   92] = 32'b01000010101100000000000000000000;
	assign	vad_gru_recurrent_weights_array[   93] = 32'b01000001110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[   94] = 32'b01000010001101000000000000000000;
	assign	vad_gru_recurrent_weights_array[   95] = 32'b11000010011011000000000000000000;
	assign	vad_gru_recurrent_weights_array[   96] = 32'b01000010100101100000000000000000;
	assign	vad_gru_recurrent_weights_array[   97] = 32'b11000010000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[   98] = 32'b01000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[   99] = 32'b01000010011001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  100] = 32'b11000010000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  101] = 32'b11000001110010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  102] = 32'b01000001010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  103] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  104] = 32'b11000010101100100000000000000000;
	assign	vad_gru_recurrent_weights_array[  105] = 32'b11000010011101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  106] = 32'b11000010100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  107] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  108] = 32'b01000001100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  109] = 32'b11000010011110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  110] = 32'b11000010100010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  111] = 32'b01000001101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  112] = 32'b11000010111000100000000000000000;
	assign	vad_gru_recurrent_weights_array[  113] = 32'b01000000101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  114] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  115] = 32'b01000010001011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  116] = 32'b11000010101100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  117] = 32'b01000001110100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  118] = 32'b11000010100111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  119] = 32'b01000001100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  120] = 32'b01000010100101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  121] = 32'b01000001101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  122] = 32'b01000001000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  123] = 32'b11000010100101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  124] = 32'b01000001101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  125] = 32'b01000010001001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  126] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  127] = 32'b11000010111011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  128] = 32'b11000001011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  129] = 32'b01000001000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  130] = 32'b01000010111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  131] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  132] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  133] = 32'b01000010000010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  134] = 32'b11000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  135] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  136] = 32'b11000011000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  137] = 32'b11000010010101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  138] = 32'b11000010010110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  139] = 32'b11000010010111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  140] = 32'b11000010111100100000000000000000;
	assign	vad_gru_recurrent_weights_array[  141] = 32'b01000010100011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  142] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  143] = 32'b11000001010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  144] = 32'b11000010100010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  145] = 32'b01000010101001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  146] = 32'b11000001110010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  147] = 32'b01000010110100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  148] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  149] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  150] = 32'b11000001101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  151] = 32'b11000001110100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  152] = 32'b01000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  153] = 32'b11000010100101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  154] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  155] = 32'b11000010111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  156] = 32'b01000001010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  157] = 32'b01000010011101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  158] = 32'b11000010100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  159] = 32'b11000010110110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  160] = 32'b11000010011111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  161] = 32'b11000010100000100000000000000000;
	assign	vad_gru_recurrent_weights_array[  162] = 32'b11000010001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  163] = 32'b11000010000011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  164] = 32'b11000010011101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  165] = 32'b11000010000111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  166] = 32'b01000010110110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  167] = 32'b11000010100101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  168] = 32'b01000010111000100000000000000000;
	assign	vad_gru_recurrent_weights_array[  169] = 32'b11000000010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  170] = 32'b01000010110110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  171] = 32'b11000001111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  172] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  173] = 32'b01000010111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  174] = 32'b01000010000111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  175] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  176] = 32'b11000011000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  177] = 32'b11000010101111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  178] = 32'b11000010110001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  179] = 32'b01000010110111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  180] = 32'b01000001000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  181] = 32'b01000001110010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  182] = 32'b01000010111001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  183] = 32'b11000010100101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  184] = 32'b11000010101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  185] = 32'b11000010010110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  186] = 32'b11000001010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  187] = 32'b11000010000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  188] = 32'b11000010000110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  189] = 32'b01000001001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  190] = 32'b01000001111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  191] = 32'b01000001001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  192] = 32'b01000010011111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  193] = 32'b01000010010011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  194] = 32'b01000010001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  195] = 32'b11000010110001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  196] = 32'b01000010100101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  197] = 32'b01000000100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  198] = 32'b01000010010010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  199] = 32'b11000011000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  200] = 32'b11000010000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  201] = 32'b11000010000011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  202] = 32'b11000001001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  203] = 32'b11000001111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  204] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  205] = 32'b11000000111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  206] = 32'b01000010100001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  207] = 32'b11000010011010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  208] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  209] = 32'b11000001101100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  210] = 32'b11000010101001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  211] = 32'b11000010011101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  212] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  213] = 32'b01000010010001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  214] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  215] = 32'b11000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  216] = 32'b01000000111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  217] = 32'b01000010011110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  218] = 32'b01000010000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  219] = 32'b11000001001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  220] = 32'b11000010000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  221] = 32'b11000010001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  222] = 32'b01000010011111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  223] = 32'b01000010111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  224] = 32'b01000010001001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  225] = 32'b01000010100000100000000000000000;
	assign	vad_gru_recurrent_weights_array[  226] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  227] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  228] = 32'b01000010011111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  229] = 32'b11000001111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  230] = 32'b11000010110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  231] = 32'b01000010100101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  232] = 32'b11000010101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  233] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  234] = 32'b01000010000110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  235] = 32'b11000001100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  236] = 32'b11000011000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  237] = 32'b01000010100010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  238] = 32'b11000000101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  239] = 32'b01000010110010100000000000000000;
	assign	vad_gru_recurrent_weights_array[  240] = 32'b11000000100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  241] = 32'b01000010101010100000000000000000;
	assign	vad_gru_recurrent_weights_array[  242] = 32'b01000010011010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  243] = 32'b01000010100111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  244] = 32'b00000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  245] = 32'b11000010011010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  246] = 32'b01000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  247] = 32'b01000010111011100000000000000000;
	assign	vad_gru_recurrent_weights_array[  248] = 32'b11000010100011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  249] = 32'b10111111100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  250] = 32'b11000010100111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  251] = 32'b11000010100010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  252] = 32'b01000010111001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  253] = 32'b11000001111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  254] = 32'b11000010101101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  255] = 32'b11000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  256] = 32'b11000010111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  257] = 32'b01000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  258] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  259] = 32'b11000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  260] = 32'b01000001001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  261] = 32'b01000010010111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  262] = 32'b11000010011011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  263] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  264] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  265] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  266] = 32'b01000010101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  267] = 32'b01000010100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  268] = 32'b01000010000011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  269] = 32'b11000010010110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  270] = 32'b01000010101111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  271] = 32'b11000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  272] = 32'b11000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  273] = 32'b01000010100111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  274] = 32'b01000001101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  275] = 32'b11000010001110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  276] = 32'b11000010011101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  277] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  278] = 32'b11000010110010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  279] = 32'b01000010110001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  280] = 32'b11000010100110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  281] = 32'b01000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  282] = 32'b11000010101011100000000000000000;
	assign	vad_gru_recurrent_weights_array[  283] = 32'b01000000101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  284] = 32'b11000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  285] = 32'b01000010010001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  286] = 32'b01000010101010100000000000000000;
	assign	vad_gru_recurrent_weights_array[  287] = 32'b01000000111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  288] = 32'b11000010100011100000000000000000;
	assign	vad_gru_recurrent_weights_array[  289] = 32'b01000010101001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  290] = 32'b01000010010101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  291] = 32'b11000010001001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  292] = 32'b01000001101100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  293] = 32'b11000001101100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  294] = 32'b11000010101110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  295] = 32'b11000010110011100000000000000000;
	assign	vad_gru_recurrent_weights_array[  296] = 32'b01000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  297] = 32'b01000010010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  298] = 32'b11000010011000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  299] = 32'b01000001011000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  300] = 32'b11000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  301] = 32'b11000010110111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  302] = 32'b01000010101010100000000000000000;
	assign	vad_gru_recurrent_weights_array[  303] = 32'b01000001100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  304] = 32'b01000010010110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  305] = 32'b01000010000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  306] = 32'b11000010111011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  307] = 32'b11000001110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  308] = 32'b01000010011101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  309] = 32'b11000010010101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  310] = 32'b01000010110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  311] = 32'b11000010100011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  312] = 32'b11000000101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  313] = 32'b11000001100010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  314] = 32'b11000010100001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  315] = 32'b11000010101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  316] = 32'b11000000111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  317] = 32'b11000010101001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  318] = 32'b11000010110101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  319] = 32'b11000010110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  320] = 32'b01000001101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  321] = 32'b11000010101001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  322] = 32'b11000010011010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  323] = 32'b01000010010010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  324] = 32'b01000001010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  325] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  326] = 32'b10111111100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  327] = 32'b11000001111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  328] = 32'b01000010000010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  329] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  330] = 32'b01000010111001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  331] = 32'b01000001100010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  332] = 32'b01000010101101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  333] = 32'b00111111100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  334] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  335] = 32'b01000010100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  336] = 32'b01000001001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  337] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  338] = 32'b11000010101000100000000000000000;
	assign	vad_gru_recurrent_weights_array[  339] = 32'b01000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  340] = 32'b01000010110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  341] = 32'b11000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  342] = 32'b01000010100110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  343] = 32'b01000001011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  344] = 32'b11000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  345] = 32'b01000010011111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  346] = 32'b11000001110110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  347] = 32'b01000001101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  348] = 32'b11000010111101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  349] = 32'b11000010110110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  350] = 32'b01000010101010100000000000000000;
	assign	vad_gru_recurrent_weights_array[  351] = 32'b11000010100111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  352] = 32'b11000001100010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  353] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  354] = 32'b11000010101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  355] = 32'b01000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  356] = 32'b11000010011101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  357] = 32'b01000001101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  358] = 32'b01000001011000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  359] = 32'b01000001100010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  360] = 32'b01000010111100100000000000000000;
	assign	vad_gru_recurrent_weights_array[  361] = 32'b01000010111101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  362] = 32'b01000001111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  363] = 32'b01000010011001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  364] = 32'b01000010111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  365] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  366] = 32'b01000010011001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  367] = 32'b01000010001010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  368] = 32'b01000010111010100000000000000000;
	assign	vad_gru_recurrent_weights_array[  369] = 32'b01000010110001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  370] = 32'b01000010100001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  371] = 32'b01000010000111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  372] = 32'b11000001101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  373] = 32'b11000010100011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  374] = 32'b01000010110010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  375] = 32'b01000000111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  376] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  377] = 32'b01000010111101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  378] = 32'b01000010001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  379] = 32'b01000001100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  380] = 32'b11000010100111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  381] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  382] = 32'b01000010101001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  383] = 32'b01000010001001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  384] = 32'b11000010110101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  385] = 32'b11000010011001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  386] = 32'b01000001110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  387] = 32'b01000010010111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  388] = 32'b01000001110110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  389] = 32'b11000010100001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  390] = 32'b11000010110111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  391] = 32'b11000010001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  392] = 32'b11000000111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  393] = 32'b11000010001011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  394] = 32'b11000010100001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  395] = 32'b01000010111100100000000000000000;
	assign	vad_gru_recurrent_weights_array[  396] = 32'b01000010001010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  397] = 32'b11000011000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  398] = 32'b11000010001101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  399] = 32'b01000010000011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  400] = 32'b01000001011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  401] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  402] = 32'b01000010000010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  403] = 32'b11000010000011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  404] = 32'b11000010000010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  405] = 32'b11000010001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  406] = 32'b11000001100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  407] = 32'b11000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  408] = 32'b01000010011111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  409] = 32'b01000010110111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  410] = 32'b01000001111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  411] = 32'b01000010111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  412] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  413] = 32'b01000001100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  414] = 32'b01000001110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  415] = 32'b11000010100011100000000000000000;
	assign	vad_gru_recurrent_weights_array[  416] = 32'b11000010000111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  417] = 32'b01000010000010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  418] = 32'b01000001001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  419] = 32'b01000001100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  420] = 32'b11000010001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  421] = 32'b01000001110110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  422] = 32'b01000001010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  423] = 32'b01000010110101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  424] = 32'b11000001001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  425] = 32'b01000010011000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  426] = 32'b11000010101001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  427] = 32'b11000010110101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  428] = 32'b11000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  429] = 32'b11000010010010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  430] = 32'b11000010010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  431] = 32'b01000010111001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  432] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  433] = 32'b11000010000010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  434] = 32'b11000010001011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  435] = 32'b11000010100010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  436] = 32'b01000001001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  437] = 32'b01000010100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  438] = 32'b01000010011001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  439] = 32'b11000010111011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  440] = 32'b11000011000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  441] = 32'b01000010000101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  442] = 32'b11000010110100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  443] = 32'b01000010100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  444] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  445] = 32'b01000000010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  446] = 32'b11000010100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  447] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  448] = 32'b11000001111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  449] = 32'b01000010101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  450] = 32'b11000010101111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  451] = 32'b11000001011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  452] = 32'b01000010010111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  453] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  454] = 32'b01000010100111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  455] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  456] = 32'b11000010011001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  457] = 32'b11000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  458] = 32'b01000010110100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  459] = 32'b11000010100010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  460] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  461] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  462] = 32'b11000010100110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  463] = 32'b01000010010011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  464] = 32'b01000010001101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  465] = 32'b01000010000001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  466] = 32'b11000010110110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  467] = 32'b01000010111001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  468] = 32'b11000001001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  469] = 32'b00111111100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  470] = 32'b01000010101111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  471] = 32'b11000010111100100000000000000000;
	assign	vad_gru_recurrent_weights_array[  472] = 32'b11000000101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  473] = 32'b11000001000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  474] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  475] = 32'b11000010111001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  476] = 32'b01000010000111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  477] = 32'b01000010100010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  478] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  479] = 32'b11000010110101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  480] = 32'b11000010010011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  481] = 32'b11000010001010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  482] = 32'b01000001110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  483] = 32'b11000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  484] = 32'b01000010010011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  485] = 32'b11000001110110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  486] = 32'b11000010001011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  487] = 32'b01000010100001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  488] = 32'b11000010001101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  489] = 32'b01000010011110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  490] = 32'b11000010110001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  491] = 32'b11000010110110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  492] = 32'b01000010100010100000000000000000;
	assign	vad_gru_recurrent_weights_array[  493] = 32'b01000010100001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  494] = 32'b00000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  495] = 32'b11000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  496] = 32'b11000011000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  497] = 32'b01000010010001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  498] = 32'b01000001111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  499] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  500] = 32'b11000010111101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  501] = 32'b01000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  502] = 32'b11000010010111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  503] = 32'b11000010100001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  504] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  505] = 32'b11000010100011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  506] = 32'b11000011000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  507] = 32'b11000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  508] = 32'b11000010100110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  509] = 32'b01000001110010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  510] = 32'b01000001100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  511] = 32'b11000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  512] = 32'b11000010110011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  513] = 32'b01000001001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  514] = 32'b11000010100101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  515] = 32'b01000010101001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  516] = 32'b01000010000110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  517] = 32'b11000000101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  518] = 32'b01000000101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  519] = 32'b01000001100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  520] = 32'b01000010000010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  521] = 32'b01000010001111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  522] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  523] = 32'b11000010101110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  524] = 32'b01000001101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  525] = 32'b01000001110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  526] = 32'b11000010110000100000000000000000;
	assign	vad_gru_recurrent_weights_array[  527] = 32'b11000001100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  528] = 32'b01000001111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  529] = 32'b01000010000111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  530] = 32'b01000010000010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  531] = 32'b11000001101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  532] = 32'b01000001101100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  533] = 32'b01000010111101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  534] = 32'b01000000111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  535] = 32'b11000010100110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  536] = 32'b11000010101000100000000000000000;
	assign	vad_gru_recurrent_weights_array[  537] = 32'b11000010001110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  538] = 32'b11000001000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  539] = 32'b00111111100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  540] = 32'b01000001101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  541] = 32'b01000010000111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  542] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  543] = 32'b11000010001011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  544] = 32'b11000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  545] = 32'b11000010010010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  546] = 32'b01000001001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  547] = 32'b11000001101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  548] = 32'b01000010011011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  549] = 32'b11000001000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  550] = 32'b11000000100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  551] = 32'b11000001010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  552] = 32'b11000001110110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  553] = 32'b01000010001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  554] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  555] = 32'b01000010010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  556] = 32'b11000010001111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  557] = 32'b01000010100011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  558] = 32'b11000010001011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  559] = 32'b01000010010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  560] = 32'b01000010110010100000000000000000;
	assign	vad_gru_recurrent_weights_array[  561] = 32'b11000010010001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  562] = 32'b01000001110110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  563] = 32'b01000010001101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  564] = 32'b01000010010001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  565] = 32'b01000010000001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  566] = 32'b11000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  567] = 32'b01000010010111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  568] = 32'b01000010111001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  569] = 32'b01000001101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  570] = 32'b10111111100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  571] = 32'b01000010100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  572] = 32'b11000001110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  573] = 32'b11000010110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  574] = 32'b01000010110100100000000000000000;
	assign	vad_gru_recurrent_weights_array[  575] = 32'b01000001110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  576] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  577] = 32'b01000010100101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  578] = 32'b11000001101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  579] = 32'b11000010110100100000000000000000;
	assign	vad_gru_recurrent_weights_array[  580] = 32'b01000001010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  581] = 32'b11000010001010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  582] = 32'b01000010001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  583] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  584] = 32'b11000001111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  585] = 32'b11000010000111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  586] = 32'b11000010101111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  587] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  588] = 32'b11000010011111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  589] = 32'b01000001001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  590] = 32'b01000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  591] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  592] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  593] = 32'b11000001011000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  594] = 32'b01000000101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  595] = 32'b01000010001010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  596] = 32'b11000010011101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  597] = 32'b11000000100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  598] = 32'b01000010010001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  599] = 32'b01000010101100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  600] = 32'b01000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  601] = 32'b11000010110101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  602] = 32'b11000001111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  603] = 32'b01000001100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  604] = 32'b11000001111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  605] = 32'b01000010001111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  606] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  607] = 32'b01000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  608] = 32'b11000010001110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  609] = 32'b11000010101100100000000000000000;
	assign	vad_gru_recurrent_weights_array[  610] = 32'b11000001100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  611] = 32'b01000010101101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  612] = 32'b11000001101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  613] = 32'b11000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  614] = 32'b01000010111011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  615] = 32'b11000001101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  616] = 32'b11000001101100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  617] = 32'b01000010000111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  618] = 32'b01000010111001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  619] = 32'b01000001001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  620] = 32'b11000010001010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  621] = 32'b01000010010110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  622] = 32'b01000010100100100000000000000000;
	assign	vad_gru_recurrent_weights_array[  623] = 32'b11000010010111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  624] = 32'b11000010100110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  625] = 32'b01000010011110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  626] = 32'b11000001110110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  627] = 32'b11000010011011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  628] = 32'b11000010110001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  629] = 32'b11000001010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  630] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  631] = 32'b11000010001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  632] = 32'b01000010011000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  633] = 32'b11000000010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  634] = 32'b11000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  635] = 32'b11000010101101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  636] = 32'b01000010100011100000000000000000;
	assign	vad_gru_recurrent_weights_array[  637] = 32'b11000010110111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  638] = 32'b01000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  639] = 32'b11000001100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  640] = 32'b01000010101001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  641] = 32'b11000001110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  642] = 32'b11000010000011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  643] = 32'b01000010110011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  644] = 32'b11000010001010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  645] = 32'b01000000111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  646] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  647] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  648] = 32'b11000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  649] = 32'b01000001100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  650] = 32'b01000010110001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  651] = 32'b11000010010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  652] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  653] = 32'b01000010110100100000000000000000;
	assign	vad_gru_recurrent_weights_array[  654] = 32'b11000010010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  655] = 32'b01000010001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  656] = 32'b11000010101001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  657] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  658] = 32'b11000010111101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  659] = 32'b01000010110110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  660] = 32'b01000000101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  661] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  662] = 32'b01000010010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  663] = 32'b01000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  664] = 32'b01000000101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  665] = 32'b11000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  666] = 32'b01000010110010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  667] = 32'b11000001100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  668] = 32'b01000001111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  669] = 32'b01000010101010100000000000000000;
	assign	vad_gru_recurrent_weights_array[  670] = 32'b11000010101100100000000000000000;
	assign	vad_gru_recurrent_weights_array[  671] = 32'b01000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  672] = 32'b01000000100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  673] = 32'b01000010001001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  674] = 32'b01000010011110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  675] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  676] = 32'b01000010011110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  677] = 32'b01000010111101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  678] = 32'b01000010101010100000000000000000;
	assign	vad_gru_recurrent_weights_array[  679] = 32'b01000010111101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  680] = 32'b11000010110101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  681] = 32'b01000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  682] = 32'b11000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  683] = 32'b01000010101110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  684] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  685] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  686] = 32'b01000010110011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  687] = 32'b01000001100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  688] = 32'b01000001100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  689] = 32'b11000010100001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  690] = 32'b01000010001001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  691] = 32'b11000010001010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  692] = 32'b01000010111001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  693] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  694] = 32'b11000010010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  695] = 32'b11000010111010100000000000000000;
	assign	vad_gru_recurrent_weights_array[  696] = 32'b11000001111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  697] = 32'b11000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  698] = 32'b11000010100100100000000000000000;
	assign	vad_gru_recurrent_weights_array[  699] = 32'b11000010110011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  700] = 32'b11000000010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  701] = 32'b11000001100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  702] = 32'b00000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  703] = 32'b01000010101100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  704] = 32'b01000010001010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  705] = 32'b01000010101011100000000000000000;
	assign	vad_gru_recurrent_weights_array[  706] = 32'b11000010111010100000000000000000;
	assign	vad_gru_recurrent_weights_array[  707] = 32'b11000001101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  708] = 32'b01000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  709] = 32'b01000010111101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  710] = 32'b01000001111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  711] = 32'b01000010011111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  712] = 32'b01000010100011100000000000000000;
	assign	vad_gru_recurrent_weights_array[  713] = 32'b01000010100001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  714] = 32'b01000010111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  715] = 32'b01000010101110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  716] = 32'b01000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  717] = 32'b11000010001011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  718] = 32'b01000010010001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  719] = 32'b01000010110011100000000000000000;
	assign	vad_gru_recurrent_weights_array[  720] = 32'b01000001111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  721] = 32'b01000010101101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  722] = 32'b11000010101101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  723] = 32'b11000001101100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  724] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  725] = 32'b01000001110100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  726] = 32'b11000001110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  727] = 32'b11000001101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  728] = 32'b01000010010011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  729] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  730] = 32'b01000010101011100000000000000000;
	assign	vad_gru_recurrent_weights_array[  731] = 32'b11000010110011100000000000000000;
	assign	vad_gru_recurrent_weights_array[  732] = 32'b11000010100010100000000000000000;
	assign	vad_gru_recurrent_weights_array[  733] = 32'b11000001001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  734] = 32'b11000010100001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  735] = 32'b11000001101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  736] = 32'b01000001101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  737] = 32'b01000010110000100000000000000000;
	assign	vad_gru_recurrent_weights_array[  738] = 32'b01000010000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  739] = 32'b01000001110010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  740] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  741] = 32'b01000001111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  742] = 32'b11000001101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  743] = 32'b11000010011111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  744] = 32'b01000001111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  745] = 32'b01000010010011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  746] = 32'b11000010111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  747] = 32'b01000001101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  748] = 32'b01000010001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  749] = 32'b11000010000111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  750] = 32'b01000010000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  751] = 32'b11000010101001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  752] = 32'b11000010100110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  753] = 32'b11000001110010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  754] = 32'b11000010010010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  755] = 32'b01000010110111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  756] = 32'b01000001011000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  757] = 32'b01000001010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  758] = 32'b11000010110110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  759] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  760] = 32'b11000010100000100000000000000000;
	assign	vad_gru_recurrent_weights_array[  761] = 32'b11000010010111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  762] = 32'b11000010101011100000000000000000;
	assign	vad_gru_recurrent_weights_array[  763] = 32'b01000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  764] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  765] = 32'b11000010000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  766] = 32'b11000010100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  767] = 32'b11000010110110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  768] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  769] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  770] = 32'b11000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  771] = 32'b11000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  772] = 32'b01000010011101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  773] = 32'b01000010111100100000000000000000;
	assign	vad_gru_recurrent_weights_array[  774] = 32'b01000010110011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  775] = 32'b11000011000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  776] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  777] = 32'b01000001100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  778] = 32'b01000010110010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  779] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  780] = 32'b11000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  781] = 32'b11000010100010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  782] = 32'b01000010100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  783] = 32'b11000010101110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  784] = 32'b11000011000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  785] = 32'b01000010001011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  786] = 32'b11000010101110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  787] = 32'b11000001100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  788] = 32'b11000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  789] = 32'b11000010110000100000000000000000;
	assign	vad_gru_recurrent_weights_array[  790] = 32'b11000010111000100000000000000000;
	assign	vad_gru_recurrent_weights_array[  791] = 32'b11000010000001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  792] = 32'b01000010101001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  793] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  794] = 32'b11000010001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  795] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  796] = 32'b11000010100101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  797] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  798] = 32'b01000001100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  799] = 32'b01000010001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  800] = 32'b01000010010010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  801] = 32'b11000010111101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  802] = 32'b01000001101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  803] = 32'b01000010111011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  804] = 32'b01000010001110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  805] = 32'b01000001100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  806] = 32'b01000001110100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  807] = 32'b11000011000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  808] = 32'b01000001001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  809] = 32'b01000000100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  810] = 32'b01000010110001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  811] = 32'b11000001011000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  812] = 32'b11000010101001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  813] = 32'b11000001010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  814] = 32'b01000001111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  815] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  816] = 32'b01000010011001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  817] = 32'b01000010100000100000000000000000;
	assign	vad_gru_recurrent_weights_array[  818] = 32'b01000010011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  819] = 32'b11000010100011100000000000000000;
	assign	vad_gru_recurrent_weights_array[  820] = 32'b01000010000011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  821] = 32'b01000010110001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  822] = 32'b01000001111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  823] = 32'b01000000111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  824] = 32'b00111111100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  825] = 32'b01000010001011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  826] = 32'b01000010101100100000000000000000;
	assign	vad_gru_recurrent_weights_array[  827] = 32'b01000010100011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  828] = 32'b01000010100101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  829] = 32'b01000010111100100000000000000000;
	assign	vad_gru_recurrent_weights_array[  830] = 32'b11000010011011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  831] = 32'b01000010101001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  832] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  833] = 32'b11000010010101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  834] = 32'b11000001100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  835] = 32'b11000010111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  836] = 32'b11000010100000100000000000000000;
	assign	vad_gru_recurrent_weights_array[  837] = 32'b01000010010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  838] = 32'b11000010010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  839] = 32'b00000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  840] = 32'b01000010101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  841] = 32'b01000010000011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  842] = 32'b01000010001101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  843] = 32'b11000010011101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  844] = 32'b01000010001110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  845] = 32'b01000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  846] = 32'b01000010110101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  847] = 32'b01000001110110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  848] = 32'b11000001110100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  849] = 32'b11000010111011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  850] = 32'b01000010101101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  851] = 32'b01000010011001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  852] = 32'b11000001001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  853] = 32'b01000000111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  854] = 32'b11000001011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  855] = 32'b00000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  856] = 32'b11000010000111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  857] = 32'b11000000100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  858] = 32'b01000001010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  859] = 32'b01000001111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  860] = 32'b10111111100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  861] = 32'b01000010111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  862] = 32'b01000010101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  863] = 32'b01000010100111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  864] = 32'b01000010111011100000000000000000;
	assign	vad_gru_recurrent_weights_array[  865] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  866] = 32'b11000010011011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  867] = 32'b01000001111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  868] = 32'b11000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  869] = 32'b11000001110010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  870] = 32'b11000010001011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  871] = 32'b01000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  872] = 32'b01000010101101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  873] = 32'b01000010100111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  874] = 32'b01000010100001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  875] = 32'b01000010110011100000000000000000;
	assign	vad_gru_recurrent_weights_array[  876] = 32'b11000010101001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  877] = 32'b01000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  878] = 32'b11000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  879] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  880] = 32'b01000001100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  881] = 32'b01000010100100100000000000000000;
	assign	vad_gru_recurrent_weights_array[  882] = 32'b00000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  883] = 32'b11000010110100100000000000000000;
	assign	vad_gru_recurrent_weights_array[  884] = 32'b01000010111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  885] = 32'b11000001100010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  886] = 32'b01000010110100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  887] = 32'b01000010110101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  888] = 32'b01000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  889] = 32'b01000010110101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  890] = 32'b01000001100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  891] = 32'b01000010011000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  892] = 32'b11000010001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  893] = 32'b01000010010111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  894] = 32'b11000010111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  895] = 32'b01000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  896] = 32'b11000010000111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  897] = 32'b11000010101001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  898] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  899] = 32'b11000010101110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  900] = 32'b11000010110001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  901] = 32'b01000010011001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  902] = 32'b11000010111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  903] = 32'b11000001101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  904] = 32'b11000010000110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  905] = 32'b01000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  906] = 32'b11000001111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  907] = 32'b11000010010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  908] = 32'b01000010110101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  909] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  910] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  911] = 32'b01000010100010100000000000000000;
	assign	vad_gru_recurrent_weights_array[  912] = 32'b01000001100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  913] = 32'b01000010110111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  914] = 32'b01000010100011100000000000000000;
	assign	vad_gru_recurrent_weights_array[  915] = 32'b01000010110100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  916] = 32'b01000010011110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  917] = 32'b11000001010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  918] = 32'b11000001101100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  919] = 32'b01000010001010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  920] = 32'b11000010000101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  921] = 32'b11000010101111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  922] = 32'b01000010000010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  923] = 32'b10111111100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  924] = 32'b11000010000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  925] = 32'b11000001010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  926] = 32'b11000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  927] = 32'b11000010001111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  928] = 32'b11000001010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  929] = 32'b01000010011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  930] = 32'b11000010100101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  931] = 32'b11000010100001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  932] = 32'b01000010011010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  933] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  934] = 32'b11000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  935] = 32'b01000010100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  936] = 32'b01000010100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  937] = 32'b11000010110101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  938] = 32'b01000010100100100000000000000000;
	assign	vad_gru_recurrent_weights_array[  939] = 32'b11000010010001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  940] = 32'b11000001111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  941] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  942] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  943] = 32'b01000001111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  944] = 32'b01000001100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  945] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  946] = 32'b11000010110111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  947] = 32'b01000010110101100000000000000000;
	assign	vad_gru_recurrent_weights_array[  948] = 32'b11000001100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  949] = 32'b11000010010101000000000000000000;
	assign	vad_gru_recurrent_weights_array[  950] = 32'b01000001101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  951] = 32'b01000010100010100000000000000000;
	assign	vad_gru_recurrent_weights_array[  952] = 32'b11000001011000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  953] = 32'b11000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  954] = 32'b01000010011011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  955] = 32'b11000010001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  956] = 32'b01000001011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  957] = 32'b01000010111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  958] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  959] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  960] = 32'b01000010001011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  961] = 32'b01000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  962] = 32'b01000001100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  963] = 32'b11000010011010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  964] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  965] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  966] = 32'b01000010001011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  967] = 32'b01000001100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  968] = 32'b01000010101001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  969] = 32'b01000010110000100000000000000000;
	assign	vad_gru_recurrent_weights_array[  970] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  971] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  972] = 32'b11000010101110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  973] = 32'b11000010001001000000000000000000;
	assign	vad_gru_recurrent_weights_array[  974] = 32'b01000010101100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  975] = 32'b00000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  976] = 32'b01000010100110100000000000000000;
	assign	vad_gru_recurrent_weights_array[  977] = 32'b11000001011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[  978] = 32'b01000010111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  979] = 32'b01000001100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  980] = 32'b11000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  981] = 32'b11000001111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  982] = 32'b11000000010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  983] = 32'b01000010101111100000000000000000;
	assign	vad_gru_recurrent_weights_array[  984] = 32'b11000010001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  985] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  986] = 32'b11000010010110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  987] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[  988] = 32'b11000010101001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  989] = 32'b11000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  990] = 32'b11000010011011000000000000000000;
	assign	vad_gru_recurrent_weights_array[  991] = 32'b01000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  992] = 32'b01000010100001100000000000000000;
	assign	vad_gru_recurrent_weights_array[  993] = 32'b11000001111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[  994] = 32'b01000000100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  995] = 32'b01000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[  996] = 32'b11000001001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  997] = 32'b01000010111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  998] = 32'b11000001111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[  999] = 32'b11000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1000] = 32'b01000010101010100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1001] = 32'b11000001101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1002] = 32'b01000010001101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1003] = 32'b01000010101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1004] = 32'b01000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1005] = 32'b11000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1006] = 32'b01000001001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1007] = 32'b01000010100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1008] = 32'b01000010000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1009] = 32'b01000010101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1010] = 32'b11000010011110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1011] = 32'b01000010100110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1012] = 32'b01000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1013] = 32'b11000010000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1014] = 32'b01000010100101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1015] = 32'b01000001111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1016] = 32'b11000010010010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1017] = 32'b01000010111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1018] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1019] = 32'b01000010111011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1020] = 32'b11000010101100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1021] = 32'b11000010010111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1022] = 32'b11000001011000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1023] = 32'b11000010000101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1024] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1025] = 32'b01000010001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1026] = 32'b11000010110110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1027] = 32'b11000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1028] = 32'b11000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1029] = 32'b01000010011001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1030] = 32'b01000010100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1031] = 32'b11000001111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1032] = 32'b11000010100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1033] = 32'b01000001111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1034] = 32'b11000010111010100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1035] = 32'b11000010101110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1036] = 32'b01000001111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1037] = 32'b11000010101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1038] = 32'b11000010001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1039] = 32'b11000010100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1040] = 32'b01000010101111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1041] = 32'b01000010011010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1042] = 32'b01000010100000100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1043] = 32'b01000010111001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1044] = 32'b01000010001001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1045] = 32'b01000010001111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1046] = 32'b01000010100011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1047] = 32'b01000010001010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1048] = 32'b11000001110100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1049] = 32'b01000010110001100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1050] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1051] = 32'b01000010011001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1052] = 32'b11000000101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1053] = 32'b01000010100101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1054] = 32'b11000001100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1055] = 32'b11000010111000100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1056] = 32'b10111111100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1057] = 32'b01000010100001100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1058] = 32'b11000001101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1059] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1060] = 32'b00111111100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1061] = 32'b11000000010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1062] = 32'b01000010000001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1063] = 32'b01000010011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1064] = 32'b11000010101001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1065] = 32'b01000010000101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1066] = 32'b11000010010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1067] = 32'b01000010101100100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1068] = 32'b01000010111001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1069] = 32'b11000010000110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1070] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1071] = 32'b11000010111001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1072] = 32'b01000010000011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1073] = 32'b01000010011010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1074] = 32'b11000000101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1075] = 32'b01000001101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1076] = 32'b11000010001110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1077] = 32'b01000010111100100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1078] = 32'b11000010111101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1079] = 32'b11000010001011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1080] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1081] = 32'b01000010111001100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1082] = 32'b01000010111101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1083] = 32'b01000010111101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1084] = 32'b11000010110010100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1085] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1086] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1087] = 32'b01000010101000100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1088] = 32'b01000010010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1089] = 32'b01000010101100100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1090] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1091] = 32'b01000010110011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1092] = 32'b01000010001010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1093] = 32'b01000010111010100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1094] = 32'b11000001000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1095] = 32'b11000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1096] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1097] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1098] = 32'b01000010110111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1099] = 32'b01000010110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1100] = 32'b01000010111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1101] = 32'b01000010100001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1102] = 32'b01000010100011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1103] = 32'b01000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1104] = 32'b01000010010111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1105] = 32'b01000010101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1106] = 32'b11000010000110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1107] = 32'b11000010011010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1108] = 32'b01000010111011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1109] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1110] = 32'b11000001100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1111] = 32'b11000010100111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1112] = 32'b01000010111101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1113] = 32'b01000001100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1114] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1115] = 32'b11000010010010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1116] = 32'b11000010000110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1117] = 32'b01000010111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1118] = 32'b11000010101010100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1119] = 32'b00111111100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1120] = 32'b01000000111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1121] = 32'b11000010011000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1122] = 32'b01000010110110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1123] = 32'b11000010100110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1124] = 32'b11000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1125] = 32'b01000001101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1126] = 32'b01000010000101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1127] = 32'b00111111100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1128] = 32'b01000001010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1129] = 32'b11000010110100100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1130] = 32'b11000010100010100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1131] = 32'b01000001111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1132] = 32'b11000010101011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1133] = 32'b01000010000001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1134] = 32'b11000010110100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1135] = 32'b11000010010011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1136] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1137] = 32'b01000010001001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1138] = 32'b01000000010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1139] = 32'b11000010111100100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1140] = 32'b01000001111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1141] = 32'b01000010100011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1142] = 32'b01000010011010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1143] = 32'b01000010101011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1144] = 32'b11000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1145] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1146] = 32'b01000010101111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1147] = 32'b11000010010111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1148] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1149] = 32'b01000010001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1150] = 32'b11000001100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1151] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1152] = 32'b11000010000001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1153] = 32'b11000010101011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1154] = 32'b11000001101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1155] = 32'b01000000111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1156] = 32'b11000010110111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1157] = 32'b11000010100010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1158] = 32'b01000001000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1159] = 32'b01000010101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1160] = 32'b11000010111011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1161] = 32'b01000010010111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1162] = 32'b11000010101001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1163] = 32'b01000010100111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1164] = 32'b11000010000101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1165] = 32'b11000001101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1166] = 32'b11000001000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1167] = 32'b11000001101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1168] = 32'b01000010010101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1169] = 32'b11000001010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1170] = 32'b01000001011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1171] = 32'b11000010001110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1172] = 32'b01000010111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1173] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1174] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1175] = 32'b01000010011000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1176] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1177] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1178] = 32'b11000000111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1179] = 32'b10111111100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1180] = 32'b01000010001101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1181] = 32'b01000001110100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1182] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1183] = 32'b01000010111100100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1184] = 32'b01000001111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1185] = 32'b01000010001111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1186] = 32'b11000010101011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1187] = 32'b01000001111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1188] = 32'b01000001001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1189] = 32'b01000010100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1190] = 32'b11000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1191] = 32'b11000000111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1192] = 32'b01000001101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1193] = 32'b01000010101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1194] = 32'b11000001010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1195] = 32'b11000010000111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1196] = 32'b11000001100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1197] = 32'b01000010101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1198] = 32'b11000010110000100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1199] = 32'b11000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1200] = 32'b11000010101010100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1201] = 32'b11000010001001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1202] = 32'b01000010010001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1203] = 32'b11000010010010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1204] = 32'b01000010111101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1205] = 32'b11000010000101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1206] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1207] = 32'b11000001111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1208] = 32'b01000001011000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1209] = 32'b01000010100111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1210] = 32'b11000010010001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1211] = 32'b11000010100000100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1212] = 32'b01000001000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1213] = 32'b11000010000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1214] = 32'b11000010000110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1215] = 32'b11000010110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1216] = 32'b01000010101010100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1217] = 32'b11000001110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1218] = 32'b11000001010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1219] = 32'b01000010000101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1220] = 32'b11000001110010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1221] = 32'b11000000101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1222] = 32'b11000010100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1223] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1224] = 32'b01000010010111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1225] = 32'b11000010011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1226] = 32'b11000001100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1227] = 32'b11000010011101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1228] = 32'b11000010011111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1229] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1230] = 32'b01000010011000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1231] = 32'b01000010100001100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1232] = 32'b01000001011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1233] = 32'b01000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1234] = 32'b01000010100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1235] = 32'b01000010111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1236] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1237] = 32'b01000010001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1238] = 32'b11000001001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1239] = 32'b01000010111001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1240] = 32'b01000001110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1241] = 32'b11000001101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1242] = 32'b01000010001110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1243] = 32'b01000010100111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1244] = 32'b11000010010101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1245] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1246] = 32'b01000010101011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1247] = 32'b01000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1248] = 32'b01000010101011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1249] = 32'b00000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1250] = 32'b01000010000110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1251] = 32'b01000010101110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1252] = 32'b01000001101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1253] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1254] = 32'b01000010111101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1255] = 32'b01000010100101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1256] = 32'b11000010100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1257] = 32'b01000001010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1258] = 32'b01000010010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1259] = 32'b01000010000001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1260] = 32'b01000010101001100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1261] = 32'b11000010010011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1262] = 32'b01000001011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1263] = 32'b11000010000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1264] = 32'b11000010010001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1265] = 32'b11000010000001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1266] = 32'b01000010111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1267] = 32'b01000010100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1268] = 32'b01000000111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1269] = 32'b01000001000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1270] = 32'b01000010100000100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1271] = 32'b01000010011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1272] = 32'b01000001101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1273] = 32'b11000001101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1274] = 32'b11000010011101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1275] = 32'b11000010010101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1276] = 32'b11000010111000100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1277] = 32'b01000010101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1278] = 32'b11000010110000100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1279] = 32'b01000010110010100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1280] = 32'b01000010000101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1281] = 32'b11000010111001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1282] = 32'b11000001110110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1283] = 32'b01000010001001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1284] = 32'b01000010100100100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1285] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1286] = 32'b11000001001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1287] = 32'b01000010011011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1288] = 32'b01000010011101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1289] = 32'b11000001011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1290] = 32'b01000010100011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1291] = 32'b11000001010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1292] = 32'b01000010101001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1293] = 32'b11000000100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1294] = 32'b01000010100010100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1295] = 32'b01000010011000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1296] = 32'b01000010101111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1297] = 32'b11000010101101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1298] = 32'b11000010010010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1299] = 32'b01000010101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1300] = 32'b11000010100101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1301] = 32'b11000010010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1302] = 32'b01000010010101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1303] = 32'b11000000111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1304] = 32'b11000010110101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1305] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1306] = 32'b01000001111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1307] = 32'b01000001111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1308] = 32'b11000001110100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1309] = 32'b11000001101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1310] = 32'b11000010011101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1311] = 32'b01000010100110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1312] = 32'b01000010101001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1313] = 32'b01000010100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1314] = 32'b11000010101101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1315] = 32'b11000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1316] = 32'b01000010111101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1317] = 32'b11000010110100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1318] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1319] = 32'b01000010111101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1320] = 32'b01000010111101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1321] = 32'b01000010111101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1322] = 32'b01000010100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1323] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1324] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1325] = 32'b11000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1326] = 32'b11000010101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1327] = 32'b01000000111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1328] = 32'b01000010001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1329] = 32'b11000010100001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1330] = 32'b11000010100000100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1331] = 32'b01000010010110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1332] = 32'b11000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1333] = 32'b01000001101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1334] = 32'b01000010110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1335] = 32'b11000010100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1336] = 32'b01000010100101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1337] = 32'b01000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1338] = 32'b11000010010101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1339] = 32'b11000001010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1340] = 32'b11000010111101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1341] = 32'b01000010000111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1342] = 32'b01000010011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1343] = 32'b11000001101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1344] = 32'b01000001100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1345] = 32'b11000001100010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1346] = 32'b11000010110000100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1347] = 32'b01000001101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1348] = 32'b11000000100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1349] = 32'b11000010010101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1350] = 32'b11000010111101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1351] = 32'b01000010000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1352] = 32'b11000001100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1353] = 32'b11000010010110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1354] = 32'b11000010101111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1355] = 32'b01000010001011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1356] = 32'b01000010100011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1357] = 32'b10111111100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1358] = 32'b11000010100001100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1359] = 32'b11000010000001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1360] = 32'b01000010001001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1361] = 32'b01000001100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1362] = 32'b01000010100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1363] = 32'b01000001111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1364] = 32'b11000010101001100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1365] = 32'b01000001111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1366] = 32'b11000010110010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1367] = 32'b11000010101101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1368] = 32'b11000001110110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1369] = 32'b01000001001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1370] = 32'b11000011000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1371] = 32'b11000010110101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1372] = 32'b01000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1373] = 32'b01000010100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1374] = 32'b11000001010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1375] = 32'b01000010001010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1376] = 32'b01000010000010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1377] = 32'b01000010111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1378] = 32'b11000001100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1379] = 32'b01000010001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1380] = 32'b01000010001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1381] = 32'b11000001000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1382] = 32'b11000001001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1383] = 32'b01000010100000100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1384] = 32'b01000010101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1385] = 32'b11000010001011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1386] = 32'b11000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1387] = 32'b01000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1388] = 32'b01000010001111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1389] = 32'b11000010000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1390] = 32'b01000001110010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1391] = 32'b01000010111101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1392] = 32'b11000001111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1393] = 32'b01000001010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1394] = 32'b01000010110010100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1395] = 32'b11000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1396] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1397] = 32'b11000001101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1398] = 32'b01000010001011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1399] = 32'b01000000111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1400] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1401] = 32'b11000001101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1402] = 32'b11000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1403] = 32'b01000010101001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1404] = 32'b11000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1405] = 32'b01000001010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1406] = 32'b11000010100100100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1407] = 32'b11000010110101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1408] = 32'b01000010111001100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1409] = 32'b01000001111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1410] = 32'b01000010111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1411] = 32'b11000001101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1412] = 32'b11000010001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1413] = 32'b11000010100011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1414] = 32'b01000010101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1415] = 32'b01000000010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1416] = 32'b01000010001111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1417] = 32'b01000010101101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1418] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1419] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1420] = 32'b11000001011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1421] = 32'b01000010101111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1422] = 32'b01000000111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1423] = 32'b01000010101110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1424] = 32'b01000000101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1425] = 32'b01000010111000100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1426] = 32'b11000010010010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1427] = 32'b01000010010110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1428] = 32'b01000001001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1429] = 32'b01000001010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1430] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1431] = 32'b01000001100010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1432] = 32'b01000010100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1433] = 32'b01000010001011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1434] = 32'b11000001101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1435] = 32'b01000000101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1436] = 32'b11000010100011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1437] = 32'b01000001101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1438] = 32'b01000001011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1439] = 32'b11000001110110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1440] = 32'b01000010110001100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1441] = 32'b01000010100010100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1442] = 32'b11000010110110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1443] = 32'b11000010111101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1444] = 32'b11000010101111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1445] = 32'b01000001100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1446] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1447] = 32'b00000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1448] = 32'b01000010111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1449] = 32'b01000010110100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1450] = 32'b01000010001101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1451] = 32'b01000010110110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1452] = 32'b11000010000010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1453] = 32'b01000010101011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1454] = 32'b01000010100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1455] = 32'b11000001011000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1456] = 32'b01000010111011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1457] = 32'b01000010001110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1458] = 32'b01000010001010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1459] = 32'b01000010110110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1460] = 32'b11000001110100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1461] = 32'b01000010101111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1462] = 32'b01000010101110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1463] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1464] = 32'b01000010011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1465] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1466] = 32'b11000010101110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1467] = 32'b11000010010110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1468] = 32'b11000010111101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1469] = 32'b01000010000010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1470] = 32'b11000010110100100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1471] = 32'b01000010011000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1472] = 32'b01000010010111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1473] = 32'b01000010110011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1474] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1475] = 32'b11000010100011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1476] = 32'b11000010010010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1477] = 32'b01000010101111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1478] = 32'b11000010100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1479] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1480] = 32'b01000010110101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1481] = 32'b01000001101010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1482] = 32'b01000010100100100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1483] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1484] = 32'b01000010011101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1485] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1486] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1487] = 32'b01000001110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1488] = 32'b11000010011110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1489] = 32'b01000010101101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1490] = 32'b01000010100100100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1491] = 32'b01000010101101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1492] = 32'b11000010001110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1493] = 32'b11000010100111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1494] = 32'b11000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1495] = 32'b01000010100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1496] = 32'b01000010111101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1497] = 32'b11000010001010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1498] = 32'b01000010010010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1499] = 32'b11000010110101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1500] = 32'b01000001100010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1501] = 32'b11000010000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1502] = 32'b11000010011110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1503] = 32'b11000010101100100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1504] = 32'b01000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1505] = 32'b00111111100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1506] = 32'b01000010101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1507] = 32'b11000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1508] = 32'b01000010111010100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1509] = 32'b01000010111011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1510] = 32'b11000010100000100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1511] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1512] = 32'b11000010101111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1513] = 32'b11000010111100100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1514] = 32'b11000010010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1515] = 32'b01000010110011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1516] = 32'b01000010100001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1517] = 32'b01000010100101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1518] = 32'b11000000010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1519] = 32'b11000010011110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1520] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1521] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1522] = 32'b11000010100101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1523] = 32'b01000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1524] = 32'b01000010100111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1525] = 32'b01000010010001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1526] = 32'b01000010001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1527] = 32'b01000010110100100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1528] = 32'b11000010100001100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1529] = 32'b11000010100011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1530] = 32'b11000010100011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1531] = 32'b01000010001011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1532] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1533] = 32'b01000010111011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1534] = 32'b11000000100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1535] = 32'b01000010100001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1536] = 32'b01000010001011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1537] = 32'b01000001101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1538] = 32'b01000010101101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1539] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1540] = 32'b01000001011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1541] = 32'b01000010011111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1542] = 32'b11000010111011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1543] = 32'b01000010111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1544] = 32'b01000010110011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1545] = 32'b01000001011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1546] = 32'b11000010110001100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1547] = 32'b01000001111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1548] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1549] = 32'b01000010100010100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1550] = 32'b01000010111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1551] = 32'b11000010001110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1552] = 32'b11000010100001100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1553] = 32'b01000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1554] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1555] = 32'b11000001111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1556] = 32'b01000001111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1557] = 32'b01000001111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1558] = 32'b11000010100010100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1559] = 32'b11000010110001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1560] = 32'b11000010001111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1561] = 32'b11000010101011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1562] = 32'b11000010100011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1563] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1564] = 32'b01000001101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1565] = 32'b11000010100100100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1566] = 32'b01000001111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1567] = 32'b11000000111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1568] = 32'b01000010101111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1569] = 32'b11000010010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1570] = 32'b11000010100000100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1571] = 32'b01000010110001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1572] = 32'b11000010001101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1573] = 32'b01000010110000100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1574] = 32'b01000010010101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1575] = 32'b01000001101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1576] = 32'b11000001000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1577] = 32'b11000001101100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1578] = 32'b11000010010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1579] = 32'b11000010001111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1580] = 32'b01000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1581] = 32'b10111111100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1582] = 32'b11000010101010100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1583] = 32'b11000001011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1584] = 32'b11000010011101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1585] = 32'b11000001011000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1586] = 32'b01000010100010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1587] = 32'b01000010110111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1588] = 32'b11000001001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1589] = 32'b11000010111100100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1590] = 32'b11000001110010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1591] = 32'b11000010000011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1592] = 32'b11000001011100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1593] = 32'b11000010101111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1594] = 32'b11000010111101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1595] = 32'b01000001110110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1596] = 32'b01000010100101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1597] = 32'b01000010010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1598] = 32'b11000010100001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1599] = 32'b11000010011000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1600] = 32'b11000010001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1601] = 32'b01000010101110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1602] = 32'b01000010110110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1603] = 32'b01000010100001100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1604] = 32'b11000010000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1605] = 32'b01000001110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1606] = 32'b01000010100011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1607] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1608] = 32'b01000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1609] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1610] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1611] = 32'b01000010010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1612] = 32'b01000001001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1613] = 32'b11000010000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1614] = 32'b01000010111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1615] = 32'b11000001010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1616] = 32'b11000001110100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1617] = 32'b11000001111000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1618] = 32'b11000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1619] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1620] = 32'b01000010110101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1621] = 32'b11000010010010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1622] = 32'b01000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1623] = 32'b01000010000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1624] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1625] = 32'b11000001010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1626] = 32'b00000000000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1627] = 32'b11000001101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1628] = 32'b01000010100110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1629] = 32'b11000010100011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1630] = 32'b11000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1631] = 32'b11000001010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1632] = 32'b11000001100010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1633] = 32'b11000010101001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1634] = 32'b01000001010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1635] = 32'b01000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1636] = 32'b01000010011001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1637] = 32'b01000010000001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1638] = 32'b01000000100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1639] = 32'b01000010100110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1640] = 32'b11000010001110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1641] = 32'b01000010100011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1642] = 32'b11000010000010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1643] = 32'b01000010100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1644] = 32'b01000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1645] = 32'b11000011000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1646] = 32'b01000010111110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1647] = 32'b11000001110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1648] = 32'b11000011000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1649] = 32'b01000010100101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1650] = 32'b11000010111100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1651] = 32'b01000010100010100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1652] = 32'b11000010001101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1653] = 32'b01000010010111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1654] = 32'b01000010000001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1655] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1656] = 32'b11000010000001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1657] = 32'b01000000100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1658] = 32'b11000010110100100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1659] = 32'b11000010001001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1660] = 32'b11000010011011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1661] = 32'b11000010101101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1662] = 32'b01000010111101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1663] = 32'b01000010001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1664] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1665] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1666] = 32'b11000010100001100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1667] = 32'b01000010010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1668] = 32'b01000001110010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1669] = 32'b11000010111110100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1670] = 32'b11000010100000100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1671] = 32'b01000010110010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1672] = 32'b11000001110010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1673] = 32'b01000010111101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1674] = 32'b01000000110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1675] = 32'b01000001001100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1676] = 32'b11000010111101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1677] = 32'b11000010101110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1678] = 32'b11000010000001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1679] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1680] = 32'b11000001100010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1681] = 32'b11000000100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1682] = 32'b01000001111010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1683] = 32'b01000010000001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1684] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1685] = 32'b01000010110000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1686] = 32'b01000000010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1687] = 32'b01000010101011100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1688] = 32'b11000010010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1689] = 32'b11000001100100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1690] = 32'b11000010100011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1691] = 32'b01000010111101100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1692] = 32'b01000010011010000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1693] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1694] = 32'b11000000010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1695] = 32'b11000010010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1696] = 32'b10111111100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1697] = 32'b11000010000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1698] = 32'b11000010001001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1699] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1700] = 32'b01000010010011000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1701] = 32'b11000010010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1702] = 32'b11000001110110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1703] = 32'b01000010001110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1704] = 32'b11000010101001100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1705] = 32'b01000010011001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1706] = 32'b01000001000100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1707] = 32'b01000010111111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1708] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1709] = 32'b01000010101111000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1710] = 32'b01000010100111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1711] = 32'b11000010000101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1712] = 32'b11000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1713] = 32'b11000010001000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1714] = 32'b01000010100001100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1715] = 32'b01000010010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1716] = 32'b01000010101001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1717] = 32'b11000010100001000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1718] = 32'b01000010111101000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1719] = 32'b11000001010100000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1720] = 32'b11000010100100100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1721] = 32'b01000010111111100000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1722] = 32'b11000001000000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1723] = 32'b11000010101000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1724] = 32'b01000010001110000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1725] = 32'b11000010010000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1726] = 32'b01000000100000000000000000000000;
	assign	vad_gru_recurrent_weights_array[ 1727] = 32'b11000010010110000000000000000000;

}
///////////////////////////////////////////////////////////////////////////////
	generate 
		genvar i, bit;
		for ( i = 0 ; i < 72 ; i = i + 1 ) 
			for ( bit = 0 ; bit < 32 ; bit = bit + 1 ) begin	
				assign vad_gru_bias[i*float+bit] = vad_gru_bias_array[i][bit];	
			end

		for ( i = 0 ; i < 1728 ; i = i + 1 ) 
			for ( bit = 0 ; bit < 32 ; bit = bit + 1 ) begin	
				assign vad_gru_input_weights[i*float+bit] = vad_gru_input_weights_array[i][bit];	
			end

		for ( i = 0 ; i < 1728 ; i = i + 1 ) 
			for ( bit = 0 ; bit < 32 ; bit = bit + 1 ) begin	
				assign vad_gru_recurrent_weights[i*float+bit] = vad_gru_recurrent_weights_array[i][bit];	
			end
	endgenerate	

	//compute update gate and reset gate  at once?



	// for compute output
	initial	begin 
		weights_scale	= 32'b0_01110111_00000000000000000000000;  // 1.f/256
		tmpsum1		= 0;
		tmpsum2		= 0;
		z 		= 0;
		r 		= 0;
		h 		= 0;
	end

	always @(posedge clk) begin
		if(index1 < N) begin

			sum 	<= vad_gru_bias[index1*float +: float];

			if(index2 < M) begin
				tmpsum1	<= vad_gru_input_weights[(index2*stride+index1)*float +: float] * dense_out[index2*float +: float];
				sum	<= tmpsum1 + sum;
				index2	<= index2 + 1;
			end

			if(index3 < M) begin
				tmpsum2	<= vad_gru_recurrent_weights[(index3*stride+index1)*float +: float] * vad_gru_state[index3*float +: float];
				sum	<= tmpsum2 + sum;
				index3	<= index3 + 1;
			end

			index1	<= index1 + 1;

			tmpz[index1*float +: float] <= weights_scale * sum;

		end
	end

	sigmoid sigforz(tmpz, z);


	always @(posedge clk) begin

		index1 =0; index2 =0; index3 = 0;

		if(index1 < N) begin

			sum <= vad_gru_bias[index1*float+N +: float];

			if(index2 < M) begin
				tmpsum1	<= vad_gru_input_weights[(N+index2*stride+index1)*float +: float] * dense_out[index2*float +: float];
				sum	<= tmpsum1 + sum;
				index2	<= index2 + 1;
			end

			if(index3 < M) begin
				tmpsum2	<= vad_gru_recurrent_weights[(N+index3*stride+index1)*float +: float] * vad_gru_state[index3*float +: float];
				sum	<= tmpsum2 + sum;
				index3	<= index3 + 1;
			end

			index1 <= index1 + 1;

			tmpr[index1*float +: float] <= weights_scale * sum;
		end
	end

	sigmoid sigforh(tmpr, r);

	integer gi;

	always @(posedge clk) begin
		gi =0; index2 =0; index3 = 0;
		
		tmpsum1 = 0; tmpsum2 = 0;
		
		if(gi < N) begin

			sum <= vad_gru_bias[2*N+gi*float+N +: float];

			if(index2 < M) begin
				tmpsum1	<= vad_gru_input_weights[(2*N+index2*stride+gi)*float +: float] * dense_out[index2*float +: float];
				sum	<= tmpsum1 + sum;
				index2	<= index2 + 1;
			end

			if(index3 < M) begin
				tmpsum2	<= vad_gru_recurrent_weights[(2*N+index3*stride+gi)*float +:32] * vad_gru_state[index3*float +: float]*r[index3*float +: float];
				sum	<= tmpsum2 + sum;
				index3	<= index3 + 1;
			end

			// tanh tanhforg1(sum, tmptmp);		// 이거 always문 안에서 모듈 선언하면 매 클럭마다 생성되니까 금지됨 듯

			h[gi*float +: float] = z[gi*float +: float]*vad_gru_state[gi*float +: float] + (one -z[gi*float +: float]) * tmptmp;

			gi <= gi + 1;
		end
	end
/*
		//always @(posedge clk) begin
	genvar gi;
	generate 
		//gi =0; index2 =0; index3 = 0;
		
		//tmpsum1 = 0; tmpsum2 = 0;
		
		if(gi < N) begin

			sum <= vad_gru_bias[2*N+gi*float+N +: float];

			if(index2 < M) begin
				tmpsum1	<= vad_gru_input_weights[(2*N+index2*stride+gi)*float +: float] * dense_out[index2*float +: float];
				sum	<= tmpsum1 + sum;
				index2	<= index2 + 1;
			end

			if(index3 < M) begin
				tmpsum2	<= vad_gru_recurrent_weights[(2*N+index3*stride+gi)*float +:32] * vad_gru_state[index3*float +: float]*r[index3*float +: float];
				sum	<= tmpsum2 + sum;
				index3	<= index3 + 1;
			end

			tanh tanhforg1(sum, tmptmp);

			h[gi*float +: float] = z[gi*float +: float]*state[gi*float +: float] + (one -z[gi*float +: float]) * tmptmp;

			gi <= gi + 1;
		end
	//end
	endgenerate
	
	assign vad_gru_state = h;

endmodule
*/
	
	assign vad_gru_state = h;

endmodule
